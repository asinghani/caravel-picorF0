//SPDX-FileCopyrightText: 2021 Anish Singhani
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0
`default_nettype none
module game_wrapper (
	VGA_R3,
	VGA_R2,
	VGA_R1,
	VGA_R0,
	VGA_G3,
	VGA_G2,
	VGA_G1,
	VGA_G0,
	VGA_B3,
	VGA_B2,
	VGA_B1,
	VGA_B0,
	VGA_VS,
	VGA_HS,
	btn_serve,
	btn_rst,
	btn0_n,
	btn1_n,
	btn2_n,
	btn3_n,
	clk_25mhz
);
	output wire VGA_R3;
	output wire VGA_R2;
	output wire VGA_R1;
	output wire VGA_R0;
	output wire VGA_G3;
	output wire VGA_G2;
	output wire VGA_G1;
	output wire VGA_G0;
	output wire VGA_B3;
	output wire VGA_B2;
	output wire VGA_B1;
	output wire VGA_B0;
	output wire VGA_VS;
	output wire VGA_HS;
	input wire btn_serve;
	input wire btn_rst;
	input wire btn0_n;
	input wire btn1_n;
	input wire btn2_n;
	input wire btn3_n;
	input wire clk_25mhz;
	wire left_up;
	wire left_down;
	wire right_up;
	wire right_down;
	wire serve;
	wire rst;
	wire [7:0] VGA_R;
	wire [7:0] VGA_G;
	wire [7:0] VGA_B;
	assign {VGA_R3, VGA_R2, VGA_R1, VGA_R0} = VGA_R[7:4];
	assign {VGA_G3, VGA_G2, VGA_G1, VGA_G0} = VGA_G[7:4];
	assign {VGA_B3, VGA_B2, VGA_B1, VGA_B0} = VGA_B[7:4];
	sync_2ff #(.WIDTH(6)) sync(
		.o_out({left_up, left_down, right_up, right_down, serve, rst}),
		.i_in({~btn0_n, ~btn1_n, ~btn2_n, ~btn3_n, btn_serve, btn_rst}),
		.i_clk(clk_25mhz),
		.i_rst('sd0)
	);
	GameTop game(
		.serve_input(serve),
		.left_move(left_up || left_down),
		.left_movedir(left_up),
		.right_move(right_up || right_down),
		.right_movedir(right_up),
		.VGA_R(VGA_R),
		.VGA_G(VGA_G),
		.VGA_B(VGA_B),
		.VGA_VS(VGA_VS),
		.VGA_HS(VGA_HS),
		.reset(rst),
		.clock(clk_25mhz)
	);
endmodule
module sync_2ff (
	o_out,
	i_in,
	i_clk,
	i_rst
);
	parameter DEFAULT = 0;
	parameter WIDTH = 1;
	output reg [WIDTH - 1:0] o_out = DEFAULT;
	input wire [WIDTH - 1:0] i_in;
	input wire i_clk;
	input wire i_rst;
	reg [WIDTH - 1:0] sync = DEFAULT;
	always @(posedge i_clk)
		if (i_rst) begin
			sync <= DEFAULT;
			o_out <= DEFAULT;
		end
		else begin
			sync <= i_in;
			o_out <= sync;
		end
endmodule
module GameTop (
	serve_input,
	left_move,
	left_movedir,
	right_move,
	right_movedir,
	VGA_R,
	VGA_G,
	VGA_B,
	VGA_VS,
	VGA_HS,
	reset,
	clock
);
	input wire serve_input;
	input wire left_move;
	input wire left_movedir;
	input wire right_move;
	input wire right_movedir;
	output wire [7:0] VGA_R;
	output wire [7:0] VGA_G;
	output wire [7:0] VGA_B;
	output wire VGA_VS;
	output wire VGA_HS;
	input wire reset;
	input wire clock;
	wire blank;
	wire [8:0] vga_row;
	wire [9:0] vga_col;
	wire [8:0] paddleLY;
	wire [8:0] paddleRY;
	wire tick_stb;
	wire [9:0] ballX;
	wire [8:0] ballY;
	wire lscored;
	wire rscored;
	wire Cnewgame;
	wire [15:0] lscore;
	wire [15:0] rscore;
	BallControl ball(
		.paddleLY(paddleLY),
		.paddleRY(paddleRY),
		.tick_stb(tick_stb),
		.serve_input(serve_input),
		.ballX(ballX),
		.ballY(ballY),
		.lscored(lscored),
		.rscored(rscored),
		.Cnewgame(Cnewgame),
		.clock(clock),
		.reset(reset)
	);
	Renderer renderer(
		.vga_r(VGA_R),
		.vga_g(VGA_G),
		.vga_b(VGA_B),
		.paddleLY(paddleLY),
		.paddleRY(paddleRY),
		.ballX(ballX),
		.ballY(ballY),
		.vga_row(vga_row),
		.vga_col(vga_col)
	);
	PaddleController left_paddle(
		.move_input(left_move),
		.movedir_input(left_movedir),
		.coord(paddleLY),
		.tick_stb(tick_stb),
		.Cnewgame(Cnewgame),
		.clock(clock)
	);
	PaddleController right_paddle(
		.move_input(right_move),
		.movedir_input(right_movedir),
		.coord(paddleRY),
		.tick_stb(tick_stb),
		.Cnewgame(Cnewgame),
		.clock(clock)
	);
	TickGen tick(
		.row(vga_row),
		.col(vga_col),
		.blank(blank),
		.tick_stb(tick_stb),
		.clock(clock)
	);
	ScoreController score(
		.lscored(lscored),
		.rscored(rscored),
		.lscore(lscore),
		.rscore(rscore),
		.Cnewgame(Cnewgame),
		.clock(clock)
	);
	vga vga(
		.HS(VGA_HS),
		.VS(VGA_VS),
		.blank(blank),
		.row(vga_row),
		.col(vga_col),
		.clock(clock),
		.reset(reset)
	);
endmodule
module vga (
	HS,
	VS,
	blank,
	row,
	col,
	clock,
	reset
);
	parameter PCLK_MULT = 1;
	output wire HS;
	output wire VS;
	output wire blank;
	output wire [8:0] row;
	output wire [9:0] col;
	input wire clock;
	input wire reset;
	wire pix_stb;
	reg [$clog2(PCLK_MULT):0] pclk_ctr;
	assign pix_stb = pclk_ctr == (PCLK_MULT - 1);
	always @(posedge clock)
		if (reset)
			pclk_ctr <= 'sd0;
		else if (pix_stb)
			pclk_ctr <= 'sd0;
		else
			pclk_ctr <= pclk_ctr + 1;
	reg [9:0] pix_ind;
	reg [9:0] line_ind;
	assign row = line_ind - 10'd31;
	assign col = pix_ind - 10'd144;
	assign HS = pix_ind >= 10'd96;
	assign VS = line_ind >= 10'd2;
	assign blank = ~(((pix_ind >= 10'd144) && (pix_ind < 10'd784)) && ((line_ind >= 10'd31) && (line_ind < 10'd511)));
	always @(posedge clock)
		if (reset) begin
			pix_ind <= 'sd0;
			line_ind <= 'sd0;
		end
		else if (pix_stb) begin
			pix_ind <= pix_ind + 1;
			if (pix_ind == 10'd799) begin
				pix_ind <= 'sd0;
				line_ind <= line_ind + 1;
				if (line_ind == 10'd520)
					line_ind <= 'sd0;
			end
		end
endmodule
module ScoreController (
	lscored,
	rscored,
	lscore,
	rscore,
	Cnewgame,
	clock
);
	input wire lscored;
	input wire rscored;
	output reg [15:0] lscore;
	output reg [15:0] rscore;
	input wire Cnewgame;
	input wire clock;
	wire [15:0] lscore_plus_one;
	wire [15:0] rscore_plus_one;
	BCDFourDigitAdd lscore_adder(
		.A(lscore),
		.B(16'h0001),
		.Sum(lscore_plus_one)
	);
	BCDFourDigitAdd rscore_adder(
		.A(rscore),
		.B(16'h0001),
		.Sum(rscore_plus_one)
	);
	always @(posedge clock)
		if (Cnewgame) begin
			lscore <= 'sd0;
			rscore <= 'sd0;
		end
		else begin
			if (lscored)
				lscore <= lscore_plus_one;
			if (rscored)
				rscore <= rscore_plus_one;
		end
endmodule
module BallControl (
	paddleLY,
	paddleRY,
	tick_stb,
	serve_input,
	ballX,
	ballY,
	lscored,
	rscored,
	Cnewgame,
	clock,
	reset
);
	input wire [8:0] paddleLY;
	input wire [8:0] paddleRY;
	input wire tick_stb;
	input wire serve_input;
	output wire [9:0] ballX;
	output wire [8:0] ballY;
	output wire lscored;
	output wire rscored;
	output wire Cnewgame;
	input wire clock;
	input wire reset;
	wire SBwall;
	wire STwall;
	wire SRpaddle;
	wire SLpaddle;
	wire Spoint;
	wire Cinplay;
	wire CVdir;
	wire CHdir;
	BallControl_cpath cpath(
		.SBwall(SBwall),
		.STwall(STwall),
		.SRpaddle(SRpaddle),
		.SLpaddle(SLpaddle),
		.Spoint(Spoint),
		.Cnewgame(Cnewgame),
		.Cinplay(Cinplay),
		.CVdir(CVdir),
		.CHdir(CHdir),
		.lscored(lscored),
		.rscored(rscored),
		.serve_input(serve_input),
		.clock(clock),
		.reset(reset)
	);
	BallControl_dpath dpath(
		.Cnewgame(Cnewgame),
		.Cinplay(Cinplay),
		.CVdir(CVdir),
		.CHdir(CHdir),
		.SBwall(SBwall),
		.STwall(STwall),
		.SRpaddle(SRpaddle),
		.SLpaddle(SLpaddle),
		.Spoint(Spoint),
		.paddleLY(paddleLY),
		.paddleRY(paddleRY),
		.tick_stb(tick_stb),
		.ballX(ballX),
		.ballY(ballY),
		.clock(clock)
	);
endmodule
module BallControl_cpath (
	SBwall,
	STwall,
	SRpaddle,
	SLpaddle,
	Spoint,
	Cnewgame,
	Cinplay,
	CVdir,
	CHdir,
	lscored,
	rscored,
	serve_input,
	clock,
	reset
);
	input wire SBwall;
	input wire STwall;
	input wire SRpaddle;
	input wire SLpaddle;
	input wire Spoint;
	output reg Cnewgame;
	output reg Cinplay;
	output reg CVdir;
	output reg CHdir;
	output reg lscored;
	output reg rscored;
	input wire serve_input;
	input wire clock;
	input wire reset;
	reg [4:0] state;
	reg [4:0] next_state;
	localparam [4:0] S_DL = 3;
	localparam [4:0] S_DR = 1;
	localparam [4:0] S_LSCORED = 7;
	localparam [4:0] S_LSCORED_WAIT = 8;
	localparam [4:0] S_RSCORED = 5;
	localparam [4:0] S_RSCORED_WAIT = 6;
	localparam [4:0] S_UL = 4;
	localparam [4:0] S_UR = 2;
	localparam [4:0] S_WAIT = 0;
	always @(*) begin
		next_state = S_WAIT;
		{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b00_0000;
		case (state)
			S_WAIT: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b10_0000;
				next_state = (serve_input ? S_DR : S_WAIT);
			end
			S_DR: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b01_1100;
				if (SRpaddle)
					next_state = S_DL;
				else if (SBwall)
					next_state = S_UR;
				else if (Spoint)
					next_state = S_LSCORED;
				else
					next_state = S_DR;
			end
			S_DL: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b01_1000;
				if (SLpaddle)
					next_state = S_DR;
				else if (SBwall)
					next_state = S_UL;
				else if (Spoint)
					next_state = S_RSCORED;
				else
					next_state = S_DL;
			end
			S_UL: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b01_0000;
				if (SLpaddle)
					next_state = S_UR;
				else if (STwall)
					next_state = S_DL;
				else if (Spoint)
					next_state = S_RSCORED;
				else
					next_state = S_UL;
			end
			S_UR: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b01_0100;
				if (SRpaddle)
					next_state = S_UL;
				else if (STwall)
					next_state = S_DR;
				else if (Spoint)
					next_state = S_LSCORED;
				else
					next_state = S_UR;
			end
			S_LSCORED: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b00_0010;
				next_state = S_LSCORED_WAIT;
			end
			S_LSCORED_WAIT: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b00_0000;
				next_state = (serve_input ? S_DR : S_LSCORED_WAIT);
			end
			S_RSCORED: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b00_0001;
				next_state = S_RSCORED_WAIT;
			end
			S_RSCORED_WAIT: begin
				{Cnewgame, Cinplay, CVdir, CHdir, lscored, rscored} = 6'b00_0000;
				next_state = (serve_input ? S_DL : S_RSCORED_WAIT);
			end
		endcase
	end
	always @(posedge clock)
		if (reset)
			state <= S_WAIT;
		else
			state <= next_state;
endmodule
module BallControl_dpath (
	Cnewgame,
	Cinplay,
	CVdir,
	CHdir,
	SBwall,
	STwall,
	SRpaddle,
	SLpaddle,
	Spoint,
	paddleLY,
	paddleRY,
	tick_stb,
	ballX,
	ballY,
	clock
);
	input wire Cnewgame;
	input wire Cinplay;
	input wire CVdir;
	input wire CHdir;
	output wire SBwall;
	output wire STwall;
	output wire SRpaddle;
	output wire SLpaddle;
	output wire Spoint;
	input wire [8:0] paddleLY;
	input wire [8:0] paddleRY;
	input wire tick_stb;
	output reg [9:0] ballX;
	output reg [8:0] ballY;
	input wire clock;
	wire is_valid_region;
	wire [9:0] nextX;
	wire [8:0] nextY;
	wire en_pos_reg;
	assign STwall = ballY < 9'd1;
	assign SBwall = ballY > ((9'd480 - 64) - 1);
	assign is_valid_region = (ballX >= 10'd1) && (ballX <= 10'd635);
	assign Spoint = ~is_valid_region;
	assign SLpaddle = ((ballX >= 60) && (ballX <= 67)) && ((ballY <= (paddleLY + 23)) && ((ballY + 63) >= paddleLY));
	assign SRpaddle = ((ballX >= 513) && (ballX <= 576)) && ((ballY <= (paddleRY + 23)) && ((ballY + 63) >= paddleRY));
	assign en_pos_reg = tick_stb || ~Cinplay;
	assign nextX = (CHdir ? ballX + 2 : ballX - 2);
	assign nextY = (CVdir ? ballY + 1 : ballY - 1);
	always @(posedge clock)
		if (en_pos_reg) begin
			ballX <= (Cinplay ? nextX : 10'd320 - 32);
			ballY <= (Cinplay ? nextY : 9'd240 - 32);
		end
endmodule
module Renderer (
	paddleLY,
	paddleRY,
	ballX,
	ballY,
	vga_row,
	vga_col,
	vga_r,
	vga_g,
	vga_b
);
	input wire [8:0] paddleLY;
	input wire [8:0] paddleRY;
	input wire [9:0] ballX;
	input wire [8:0] ballY;
	input wire [8:0] vga_row;
	input wire [9:0] vga_col;
	output reg [7:0] vga_r;
	output reg [7:0] vga_g;
	output reg [7:0] vga_b;
	wire ispaddleL;
	wire ispaddleR;
	wire isball;
	assign ispaddleL = (((vga_row >= paddleLY) && (vga_row <= (paddleLY + 23))) && (vga_col >= 60)) && (vga_col <= 67);
	assign ispaddleR = (((vga_row >= paddleRY) && (vga_row <= (paddleRY + 23))) && (vga_col >= 577)) && (vga_col <= 584);
	assign isball = (((vga_row >= ballY) && (vga_row <= (ballY + 63))) && (vga_col >= ballX)) && (vga_col <= (ballX + 63));
	wire [23:0] ballrom_out;
	BallROM ball(
		.col(vga_col - ballX),
		.row(vga_row - ballY),
		.color(ballrom_out)
	);
	always @(*)
		if (isball)
			{vga_r, vga_g, vga_b} = ballrom_out;
		else if (ispaddleL)
			{vga_r, vga_g, vga_b} = 24'h00FFFF;
		else if (ispaddleR)
			{vga_r, vga_g, vga_b} = 24'h00FFFF;
		else
			{vga_r, vga_g, vga_b} = 24'h000000;
endmodule
module PaddleController (
	move_input,
	movedir_input,
	coord,
	tick_stb,
	Cnewgame,
	clock
);
	input wire move_input;
	input wire movedir_input;
	output reg [8:0] coord;
	input wire tick_stb;
	input wire Cnewgame;
	input wire clock;
	wire [8:0] next_coord;
	assign next_coord = (movedir_input ? coord - 5 : coord + 5);
	always @(posedge clock)
		if (Cnewgame)
			coord <= 'sd0;
		else if ((tick_stb && move_input) && (next_coord <= 456))
			coord <= next_coord;
endmodule
module TickGen (
	row,
	col,
	blank,
	tick_stb,
	clock
);
	input wire [8:0] row;
	input wire [9:0] col;
	input wire blank;
	output wire tick_stb;
	input wire clock;
	assign tick_stb = ((row == 9'd479) && (col == 10'd639)) && !blank;
endmodule
module BCDFourDigitAdd (
	A,
	B,
	Sum
);
	input wire [15:0] A;
	input wire [15:0] B;
	output wire [15:0] Sum;
	wire [2:0] carry;
	BCDOneDigitAdd add0(
		.A(A[3:0]),
		.B(B[3:0]),
		.Sum(Sum[3:0]),
		.Cin('sd0),
		.Cout(carry[0])
	);
	BCDOneDigitAdd add1(
		.A(A[7:4]),
		.B(B[7:4]),
		.Sum(Sum[7:4]),
		.Cin(carry[0]),
		.Cout(carry[1])
	);
	BCDOneDigitAdd add2(
		.A(A[11:8]),
		.B(B[11:8]),
		.Sum(Sum[11:8]),
		.Cin(carry[1]),
		.Cout(carry[2])
	);
	BCDOneDigitAdd add3(
		.A(A[15:12]),
		.B(B[15:12]),
		.Sum(Sum[15:12]),
		.Cin(carry[2]),
		.Cout()
	);
endmodule
module BCDOneDigitAdd (
	A,
	B,
	Cin,
	Sum,
	Cout
);
	input wire [3:0] A;
	input wire [3:0] B;
	input wire Cin;
	output wire [3:0] Sum;
	output wire Cout;
	wire [4:0] bin_sum;
	assign bin_sum = (A + B) + Cin;
	assign Cout = bin_sum >= 5'd10;
	assign Sum = (Cout ? bin_sum - 5'd10 : bin_sum);
endmodule
module BallROM (
	col,
	row,
	color
);
	input wire [5:0] col;
	input wire [5:0] row;
	output reg [23:0] color;
	always @(*)
		case ({col, row})
			{6'd0, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd0}: color = {8'd64, 8'd64, 8'd64};
			{6'd27, 6'd0}: color = {8'd64, 8'd64, 8'd64};
			{6'd28, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd29, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd30, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd31, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd32, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd33, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd34, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd35, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd36, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd37, 6'd0}: color = {8'd128, 8'd128, 8'd128};
			{6'd38, 6'd0}: color = {8'd64, 8'd64, 8'd64};
			{6'd39, 6'd0}: color = {8'd64, 8'd64, 8'd64};
			{6'd40, 6'd0}: color = {8'd64, 8'd64, 8'd64};
			{6'd41, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd0}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd1}: color = {8'd64, 8'd64, 8'd64};
			{6'd23, 6'd1}: color = {8'd64, 8'd64, 8'd64};
			{6'd24, 6'd1}: color = {8'd128, 8'd128, 8'd128};
			{6'd25, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd32, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd33, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd34, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd39, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd40, 6'd1}: color = {8'd192, 8'd192, 8'd192};
			{6'd41, 6'd1}: color = {8'd128, 8'd128, 8'd128};
			{6'd42, 6'd1}: color = {8'd128, 8'd128, 8'd128};
			{6'd43, 6'd1}: color = {8'd64, 8'd64, 8'd64};
			{6'd44, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd1}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd2}: color = {8'd64, 8'd64, 8'd64};
			{6'd21, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd22, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd31, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd32, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd33, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd34, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd35, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd36, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd39, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd40, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd41, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd42, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd43, 6'd2}: color = {8'd192, 8'd192, 8'd192};
			{6'd44, 6'd2}: color = {8'd128, 8'd128, 8'd128};
			{6'd45, 6'd2}: color = {8'd64, 8'd64, 8'd64};
			{6'd46, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd2}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd19, 6'd3}: color = {8'd128, 8'd128, 8'd128};
			{6'd20, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd3}: color = {8'd128, 8'd128, 8'd128};
			{6'd26, 6'd3}: color = {8'd128, 8'd128, 8'd128};
			{6'd27, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd28, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd29, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd30, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd31, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd32, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd33, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd34, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd35, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd36, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd37, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd38, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd39, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd40, 6'd3}: color = {8'd128, 8'd128, 8'd128};
			{6'd41, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd42, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd43, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd44, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd45, 6'd3}: color = {8'd192, 8'd192, 8'd192};
			{6'd46, 6'd3}: color = {8'd128, 8'd128, 8'd128};
			{6'd47, 6'd3}: color = {8'd64, 8'd64, 8'd64};
			{6'd48, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd3}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd4}: color = {8'd64, 8'd64, 8'd64};
			{6'd17, 6'd4}: color = {8'd128, 8'd128, 8'd128};
			{6'd18, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd4}: color = {8'd128, 8'd128, 8'd128};
			{6'd23, 6'd4}: color = {8'd64, 8'd64, 8'd64};
			{6'd24, 6'd4}: color = {8'd64, 8'd64, 8'd64};
			{6'd25, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd27, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd28, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd29, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd30, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd31, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd32, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd33, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd34, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd35, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd36, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd37, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd38, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd39, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd40, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd4}: color = {8'd64, 8'd64, 8'd64};
			{6'd42, 6'd4}: color = {8'd64, 8'd64, 8'd64};
			{6'd43, 6'd4}: color = {8'd128, 8'd128, 8'd128};
			{6'd44, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd45, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd46, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd47, 6'd4}: color = {8'd192, 8'd192, 8'd192};
			{6'd48, 6'd4}: color = {8'd128, 8'd128, 8'd128};
			{6'd49, 6'd4}: color = {8'd64, 8'd64, 8'd64};
			{6'd50, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd4}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd5}: color = {8'd128, 8'd128, 8'd128};
			{6'd16, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd5}: color = {8'd128, 8'd128, 8'd128};
			{6'd21, 6'd5}: color = {8'd64, 8'd64, 8'd64};
			{6'd22, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd5}: color = {8'd128, 8'd128, 8'd64};
			{6'd27, 6'd5}: color = {8'd192, 8'd128, 8'd64};
			{6'd28, 6'd5}: color = {8'd192, 8'd128, 8'd64};
			{6'd29, 6'd5}: color = {8'd128, 8'd128, 8'd64};
			{6'd30, 6'd5}: color = {8'd128, 8'd128, 8'd64};
			{6'd31, 6'd5}: color = {8'd64, 8'd64, 8'd64};
			{6'd32, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd33, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd34, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd35, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd36, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd37, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd38, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd39, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd40, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd5}: color = {8'd64, 8'd64, 8'd64};
			{6'd45, 6'd5}: color = {8'd128, 8'd128, 8'd128};
			{6'd46, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd47, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd48, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd49, 6'd5}: color = {8'd192, 8'd192, 8'd192};
			{6'd50, 6'd5}: color = {8'd128, 8'd128, 8'd128};
			{6'd51, 6'd5}: color = {8'd64, 8'd64, 8'd64};
			{6'd52, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd5}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd6}: color = {8'd64, 8'd64, 8'd64};
			{6'd14, 6'd6}: color = {8'd128, 8'd128, 8'd128};
			{6'd15, 6'd6}: color = {8'd192, 8'd192, 8'd192};
			{6'd16, 6'd6}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd6}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd6}: color = {8'd128, 8'd128, 8'd128};
			{6'd19, 6'd6}: color = {8'd64, 8'd64, 8'd64};
			{6'd20, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd6}: color = {8'd64, 8'd64, 8'd64};
			{6'd26, 6'd6}: color = {8'd128, 8'd128, 8'd128};
			{6'd27, 6'd6}: color = {8'd64, 8'd64, 8'd64};
			{6'd28, 6'd6}: color = {8'd128, 8'd128, 8'd64};
			{6'd29, 6'd6}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd6}: color = {8'd128, 8'd128, 8'd64};
			{6'd31, 6'd6}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd6}: color = {8'd128, 8'd128, 8'd64};
			{6'd33, 6'd6}: color = {8'd128, 8'd128, 8'd64};
			{6'd34, 6'd6}: color = {8'd64, 8'd64, 8'd64};
			{6'd35, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd36, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd37, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd38, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd39, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd40, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd6}: color = {8'd64, 8'd64, 8'd64};
			{6'd47, 6'd6}: color = {8'd128, 8'd128, 8'd128};
			{6'd48, 6'd6}: color = {8'd192, 8'd192, 8'd192};
			{6'd49, 6'd6}: color = {8'd192, 8'd192, 8'd192};
			{6'd50, 6'd6}: color = {8'd192, 8'd192, 8'd192};
			{6'd51, 6'd6}: color = {8'd192, 8'd192, 8'd192};
			{6'd52, 6'd6}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd6}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd7}: color = {8'd64, 8'd64, 8'd64};
			{6'd13, 6'd7}: color = {8'd192, 8'd192, 8'd192};
			{6'd14, 6'd7}: color = {8'd192, 8'd192, 8'd192};
			{6'd15, 6'd7}: color = {8'd192, 8'd192, 8'd192};
			{6'd16, 6'd7}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd7}: color = {8'd64, 8'd64, 8'd64};
			{6'd18, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd27, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd28, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd29, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd30, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd31, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd32, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd33, 6'd7}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd7}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd7}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd7}: color = {8'd128, 8'd128, 8'd64};
			{6'd37, 6'd7}: color = {8'd64, 8'd64, 8'd64};
			{6'd38, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd39, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd40, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd7}: color = {8'd64, 8'd64, 8'd64};
			{6'd49, 6'd7}: color = {8'd128, 8'd128, 8'd128};
			{6'd50, 6'd7}: color = {8'd192, 8'd192, 8'd192};
			{6'd51, 6'd7}: color = {8'd192, 8'd192, 8'd192};
			{6'd52, 6'd7}: color = {8'd192, 8'd192, 8'd192};
			{6'd53, 6'd7}: color = {8'd128, 8'd128, 8'd128};
			{6'd54, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd7}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd8}: color = {8'd64, 8'd64, 8'd64};
			{6'd12, 6'd8}: color = {8'd192, 8'd192, 8'd192};
			{6'd13, 6'd8}: color = {8'd192, 8'd192, 8'd192};
			{6'd14, 6'd8}: color = {8'd192, 8'd192, 8'd192};
			{6'd15, 6'd8}: color = {8'd128, 8'd128, 8'd128};
			{6'd16, 6'd8}: color = {8'd64, 8'd64, 8'd64};
			{6'd17, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd8}: color = {8'd128, 8'd128, 8'd64};
			{6'd26, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd27, 6'd8}: color = {8'd128, 8'd64, 8'd0};
			{6'd28, 6'd8}: color = {8'd128, 8'd128, 8'd64};
			{6'd29, 6'd8}: color = {8'd128, 8'd128, 8'd64};
			{6'd30, 6'd8}: color = {8'd128, 8'd128, 8'd64};
			{6'd31, 6'd8}: color = {8'd128, 8'd128, 8'd64};
			{6'd32, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd33, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd38, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd39, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd40, 6'd8}: color = {8'd192, 8'd128, 8'd64};
			{6'd41, 6'd8}: color = {8'd192, 8'd128, 8'd128};
			{6'd42, 6'd8}: color = {8'd128, 8'd128, 8'd64};
			{6'd43, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd8}: color = {8'd128, 8'd128, 8'd128};
			{6'd51, 6'd8}: color = {8'd192, 8'd192, 8'd192};
			{6'd52, 6'd8}: color = {8'd192, 8'd192, 8'd192};
			{6'd53, 6'd8}: color = {8'd192, 8'd192, 8'd192};
			{6'd54, 6'd8}: color = {8'd128, 8'd128, 8'd128};
			{6'd55, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd8}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd9}: color = {8'd128, 8'd128, 8'd128};
			{6'd11, 6'd9}: color = {8'd192, 8'd192, 8'd192};
			{6'd12, 6'd9}: color = {8'd192, 8'd192, 8'd192};
			{6'd13, 6'd9}: color = {8'd192, 8'd192, 8'd192};
			{6'd14, 6'd9}: color = {8'd128, 8'd128, 8'd128};
			{6'd15, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd9}: color = {8'd64, 8'd64, 8'd64};
			{6'd25, 6'd9}: color = {8'd128, 8'd128, 8'd128};
			{6'd26, 6'd9}: color = {8'd128, 8'd128, 8'd64};
			{6'd27, 6'd9}: color = {8'd128, 8'd128, 8'd64};
			{6'd28, 6'd9}: color = {8'd128, 8'd128, 8'd64};
			{6'd29, 6'd9}: color = {8'd128, 8'd64, 8'd64};
			{6'd30, 6'd9}: color = {8'd128, 8'd64, 8'd64};
			{6'd31, 6'd9}: color = {8'd128, 8'd64, 8'd64};
			{6'd32, 6'd9}: color = {8'd128, 8'd128, 8'd64};
			{6'd33, 6'd9}: color = {8'd128, 8'd128, 8'd64};
			{6'd34, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd38, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd39, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd40, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd41, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd42, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd43, 6'd9}: color = {8'd192, 8'd128, 8'd64};
			{6'd44, 6'd9}: color = {8'd64, 8'd64, 8'd64};
			{6'd45, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd9}: color = {8'd64, 8'd64, 8'd64};
			{6'd52, 6'd9}: color = {8'd192, 8'd192, 8'd192};
			{6'd53, 6'd9}: color = {8'd192, 8'd192, 8'd192};
			{6'd54, 6'd9}: color = {8'd192, 8'd192, 8'd192};
			{6'd55, 6'd9}: color = {8'd128, 8'd128, 8'd128};
			{6'd56, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd9}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd10}: color = {8'd64, 8'd64, 8'd64};
			{6'd10, 6'd10}: color = {8'd192, 8'd192, 8'd192};
			{6'd11, 6'd10}: color = {8'd192, 8'd192, 8'd192};
			{6'd12, 6'd10}: color = {8'd192, 8'd192, 8'd192};
			{6'd13, 6'd10}: color = {8'd64, 8'd64, 8'd64};
			{6'd14, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd10}: color = {8'd64, 8'd64, 8'd0};
			{6'd25, 6'd10}: color = {8'd192, 8'd128, 8'd128};
			{6'd26, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd27, 6'd10}: color = {8'd128, 8'd64, 8'd64};
			{6'd28, 6'd10}: color = {8'd128, 8'd64, 8'd64};
			{6'd29, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd30, 6'd10}: color = {8'd128, 8'd64, 8'd64};
			{6'd31, 6'd10}: color = {8'd128, 8'd64, 8'd64};
			{6'd32, 6'd10}: color = {8'd64, 8'd64, 8'd64};
			{6'd33, 6'd10}: color = {8'd128, 8'd64, 8'd64};
			{6'd34, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd35, 6'd10}: color = {8'd128, 8'd64, 8'd64};
			{6'd36, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd37, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd38, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd39, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd40, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd41, 6'd10}: color = {8'd192, 8'd128, 8'd64};
			{6'd42, 6'd10}: color = {8'd192, 8'd128, 8'd64};
			{6'd43, 6'd10}: color = {8'd192, 8'd128, 8'd64};
			{6'd44, 6'd10}: color = {8'd192, 8'd128, 8'd64};
			{6'd45, 6'd10}: color = {8'd128, 8'd128, 8'd64};
			{6'd46, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd10}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd10}: color = {8'd192, 8'd192, 8'd192};
			{6'd54, 6'd10}: color = {8'd192, 8'd192, 8'd192};
			{6'd55, 6'd10}: color = {8'd192, 8'd192, 8'd192};
			{6'd56, 6'd10}: color = {8'd128, 8'd128, 8'd128};
			{6'd57, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd10}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd11}: color = {8'd64, 8'd64, 8'd64};
			{6'd9, 6'd11}: color = {8'd192, 8'd192, 8'd192};
			{6'd10, 6'd11}: color = {8'd192, 8'd192, 8'd192};
			{6'd11, 6'd11}: color = {8'd192, 8'd192, 8'd192};
			{6'd12, 6'd11}: color = {8'd64, 8'd64, 8'd64};
			{6'd13, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd11}: color = {8'd64, 8'd64, 8'd64};
			{6'd25, 6'd11}: color = {8'd64, 8'd64, 8'd64};
			{6'd26, 6'd11}: color = {8'd64, 8'd64, 8'd64};
			{6'd27, 6'd11}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd11}: color = {8'd192, 8'd128, 8'd128};
			{6'd29, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd30, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd31, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd32, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd33, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd34, 6'd11}: color = {8'd128, 8'd64, 8'd64};
			{6'd35, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd36, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd37, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd38, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd39, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd40, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd41, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd42, 6'd11}: color = {8'd192, 8'd128, 8'd64};
			{6'd43, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd44, 6'd11}: color = {8'd128, 8'd128, 8'd0};
			{6'd45, 6'd11}: color = {8'd192, 8'd128, 8'd64};
			{6'd46, 6'd11}: color = {8'd128, 8'd128, 8'd64};
			{6'd47, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd11}: color = {8'd64, 8'd64, 8'd64};
			{6'd54, 6'd11}: color = {8'd192, 8'd192, 8'd192};
			{6'd55, 6'd11}: color = {8'd192, 8'd192, 8'd192};
			{6'd56, 6'd11}: color = {8'd192, 8'd192, 8'd192};
			{6'd57, 6'd11}: color = {8'd128, 8'd128, 8'd128};
			{6'd58, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd11}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd12}: color = {8'd64, 8'd64, 8'd64};
			{6'd8, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd10, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd11, 6'd12}: color = {8'd64, 8'd64, 8'd64};
			{6'd12, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd12}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd12}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd12}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd12}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd12}: color = {8'd192, 8'd128, 8'd0};
			{6'd33, 6'd12}: color = {8'd128, 8'd128, 8'd0};
			{6'd34, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd35, 6'd12}: color = {8'd64, 8'd64, 8'd0};
			{6'd36, 6'd12}: color = {8'd64, 8'd64, 8'd0};
			{6'd37, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd38, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd39, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd40, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd41, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd42, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd43, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd44, 6'd12}: color = {8'd128, 8'd64, 8'd64};
			{6'd45, 6'd12}: color = {8'd128, 8'd64, 8'd0};
			{6'd46, 6'd12}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd12}: color = {8'd128, 8'd128, 8'd64};
			{6'd48, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd12}: color = {8'd64, 8'd64, 8'd64};
			{6'd55, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd56, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd57, 6'd12}: color = {8'd192, 8'd192, 8'd192};
			{6'd58, 6'd12}: color = {8'd64, 8'd64, 8'd64};
			{6'd59, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd12}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd13}: color = {8'd128, 8'd128, 8'd128};
			{6'd8, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd10, 6'd13}: color = {8'd128, 8'd128, 8'd128};
			{6'd11, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd13}: color = {8'd128, 8'd128, 8'd128};
			{6'd26, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd13}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd13}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd13}: color = {8'd192, 8'd128, 8'd128};
			{6'd33, 6'd13}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd13}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd13}: color = {8'd128, 8'd128, 8'd64};
			{6'd36, 6'd13}: color = {8'd128, 8'd64, 8'd0};
			{6'd37, 6'd13}: color = {8'd128, 8'd64, 8'd0};
			{6'd38, 6'd13}: color = {8'd128, 8'd64, 8'd0};
			{6'd39, 6'd13}: color = {8'd128, 8'd64, 8'd64};
			{6'd40, 6'd13}: color = {8'd128, 8'd64, 8'd64};
			{6'd41, 6'd13}: color = {8'd128, 8'd64, 8'd64};
			{6'd42, 6'd13}: color = {8'd128, 8'd128, 8'd64};
			{6'd43, 6'd13}: color = {8'd128, 8'd128, 8'd64};
			{6'd44, 6'd13}: color = {8'd64, 8'd64, 8'd0};
			{6'd45, 6'd13}: color = {8'd64, 8'd64, 8'd0};
			{6'd46, 6'd13}: color = {8'd128, 8'd128, 8'd0};
			{6'd47, 6'd13}: color = {8'd192, 8'd128, 8'd128};
			{6'd48, 6'd13}: color = {8'd64, 8'd64, 8'd64};
			{6'd49, 6'd13}: color = {8'd128, 8'd64, 8'd64};
			{6'd50, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd13}: color = {8'd64, 8'd64, 8'd64};
			{6'd56, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd57, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd58, 6'd13}: color = {8'd192, 8'd192, 8'd192};
			{6'd59, 6'd13}: color = {8'd64, 8'd64, 8'd64};
			{6'd60, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd13}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd14}: color = {8'd128, 8'd128, 8'd128};
			{6'd7, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd8, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd14}: color = {8'd128, 8'd128, 8'd128};
			{6'd10, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd14}: color = {8'd128, 8'd128, 8'd128};
			{6'd25, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd32, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd14}: color = {8'd192, 8'd128, 8'd128};
			{6'd42, 6'd14}: color = {8'd192, 8'd128, 8'd128};
			{6'd43, 6'd14}: color = {8'd64, 8'd64, 8'd64};
			{6'd44, 6'd14}: color = {8'd128, 8'd64, 8'd64};
			{6'd45, 6'd14}: color = {8'd192, 8'd128, 8'd128};
			{6'd46, 6'd14}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd14}: color = {8'd192, 8'd128, 8'd64};
			{6'd48, 6'd14}: color = {8'd128, 8'd64, 8'd64};
			{6'd49, 6'd14}: color = {8'd192, 8'd192, 8'd128};
			{6'd50, 6'd14}: color = {8'd128, 8'd128, 8'd64};
			{6'd51, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd14}: color = {8'd128, 8'd128, 8'd128};
			{6'd57, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd58, 6'd14}: color = {8'd192, 8'd192, 8'd192};
			{6'd59, 6'd14}: color = {8'd128, 8'd128, 8'd128};
			{6'd60, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd14}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd15}: color = {8'd64, 8'd64, 8'd64};
			{6'd6, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd8, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd15}: color = {8'd64, 8'd64, 8'd64};
			{6'd10, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd34, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd15}: color = {8'd192, 8'd128, 8'd128};
			{6'd42, 6'd15}: color = {8'd128, 8'd64, 8'd64};
			{6'd43, 6'd15}: color = {8'd128, 8'd128, 8'd64};
			{6'd44, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd15}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd15}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd15}: color = {8'd128, 8'd128, 8'd64};
			{6'd48, 6'd15}: color = {8'd192, 8'd128, 8'd64};
			{6'd49, 6'd15}: color = {8'd128, 8'd128, 8'd64};
			{6'd50, 6'd15}: color = {8'd128, 8'd128, 8'd64};
			{6'd51, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd15}: color = {8'd128, 8'd128, 8'd128};
			{6'd58, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd59, 6'd15}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd15}: color = {8'd64, 8'd64, 8'd64};
			{6'd61, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd15}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd16}: color = {8'd128, 8'd128, 8'd128};
			{6'd6, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd8, 6'd16}: color = {8'd64, 8'd64, 8'd64};
			{6'd9, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd16}: color = {8'd192, 8'd128, 8'd128};
			{6'd42, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd44, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd16}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd16}: color = {8'd192, 8'd128, 8'd128};
			{6'd47, 6'd16}: color = {8'd128, 8'd64, 8'd0};
			{6'd48, 6'd16}: color = {8'd128, 8'd128, 8'd64};
			{6'd49, 6'd16}: color = {8'd192, 8'd128, 8'd64};
			{6'd50, 6'd16}: color = {8'd192, 8'd128, 8'd64};
			{6'd51, 6'd16}: color = {8'd128, 8'd64, 8'd64};
			{6'd52, 6'd16}: color = {8'd0, 8'd64, 8'd0};
			{6'd53, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd16}: color = {8'd64, 8'd64, 8'd64};
			{6'd58, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd59, 6'd16}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd16}: color = {8'd128, 8'd128, 8'd128};
			{6'd61, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd16}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd17}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd17}: color = {8'd128, 8'd128, 8'd128};
			{6'd8, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd17}: color = {8'd64, 8'd64, 8'd64};
			{6'd23, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd42, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd43, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd17}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd17}: color = {8'd128, 8'd128, 8'd128};
			{6'd47, 6'd17}: color = {8'd128, 8'd64, 8'd0};
			{6'd48, 6'd17}: color = {8'd128, 8'd128, 8'd64};
			{6'd49, 6'd17}: color = {8'd128, 8'd128, 8'd64};
			{6'd50, 6'd17}: color = {8'd192, 8'd128, 8'd64};
			{6'd51, 6'd17}: color = {8'd128, 8'd128, 8'd64};
			{6'd52, 6'd17}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd17}: color = {8'd128, 8'd128, 8'd128};
			{6'd59, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd17}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd17}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd17}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd18}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd18}: color = {8'd64, 8'd64, 8'd64};
			{6'd8, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd26, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd33, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd18}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd18}: color = {8'd192, 8'd128, 8'd128};
			{6'd47, 6'd18}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd18}: color = {8'd128, 8'd128, 8'd0};
			{6'd49, 6'd18}: color = {8'd128, 8'd128, 8'd64};
			{6'd50, 6'd18}: color = {8'd192, 8'd128, 8'd64};
			{6'd51, 6'd18}: color = {8'd192, 8'd128, 8'd64};
			{6'd52, 6'd18}: color = {8'd64, 8'd64, 8'd0};
			{6'd53, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd18}: color = {8'd64, 8'd64, 8'd64};
			{6'd59, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd18}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd18}: color = {8'd128, 8'd128, 8'd128};
			{6'd62, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd18}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd19}: color = {8'd64, 8'd64, 8'd64};
			{6'd4, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd19}: color = {8'd128, 8'd128, 8'd128};
			{6'd7, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd32, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd33, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd19}: color = {8'd192, 8'd192, 8'd128};
			{6'd47, 6'd19}: color = {8'd128, 8'd64, 8'd64};
			{6'd48, 6'd19}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd19}: color = {8'd128, 8'd64, 8'd0};
			{6'd50, 6'd19}: color = {8'd192, 8'd128, 8'd64};
			{6'd51, 6'd19}: color = {8'd192, 8'd128, 8'd64};
			{6'd52, 6'd19}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd19}: color = {8'd128, 8'd128, 8'd128};
			{6'd60, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd19}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd19}: color = {8'd64, 8'd64, 8'd64};
			{6'd63, 6'd19}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd20}: color = {8'd128, 8'd128, 8'd128};
			{6'd4, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd20}: color = {8'd64, 8'd64, 8'd64};
			{6'd7, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd20}: color = {8'd64, 8'd64, 8'd64};
			{6'd22, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd32, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd20}: color = {8'd192, 8'd192, 8'd128};
			{6'd47, 6'd20}: color = {8'd128, 8'd128, 8'd64};
			{6'd48, 6'd20}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd20}: color = {8'd128, 8'd64, 8'd0};
			{6'd50, 6'd20}: color = {8'd192, 8'd128, 8'd64};
			{6'd51, 6'd20}: color = {8'd192, 8'd128, 8'd64};
			{6'd52, 6'd20}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd20}: color = {8'd64, 8'd64, 8'd64};
			{6'd60, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd20}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd20}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd20}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd21}: color = {8'd128, 8'd128, 8'd128};
			{6'd6, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd21}: color = {8'd64, 8'd64, 8'd64};
			{6'd22, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd44, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd21}: color = {8'd192, 8'd192, 8'd128};
			{6'd47, 6'd21}: color = {8'd128, 8'd64, 8'd64};
			{6'd48, 6'd21}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd21}: color = {8'd128, 8'd64, 8'd0};
			{6'd50, 6'd21}: color = {8'd192, 8'd128, 8'd64};
			{6'd51, 6'd21}: color = {8'd128, 8'd128, 8'd64};
			{6'd52, 6'd21}: color = {8'd64, 8'd64, 8'd0};
			{6'd53, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd21}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd21}: color = {8'd128, 8'd128, 8'd128};
			{6'd61, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd21}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd21}: color = {8'd64, 8'd64, 8'd64};
			{6'd0, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd22}: color = {8'd64, 8'd64, 8'd64};
			{6'd3, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd22}: color = {8'd128, 8'd128, 8'd128};
			{6'd6, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd22}: color = {8'd128, 8'd128, 8'd128};
			{6'd22, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd24, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd26, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd44, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd22}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd22}: color = {8'd192, 8'd128, 8'd128};
			{6'd47, 6'd22}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd22}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd22}: color = {8'd64, 8'd64, 8'd0};
			{6'd50, 6'd22}: color = {8'd128, 8'd128, 8'd64};
			{6'd51, 6'd22}: color = {8'd128, 8'd128, 8'd64};
			{6'd52, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd22}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd22}: color = {8'd64, 8'd64, 8'd64};
			{6'd61, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd22}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd22}: color = {8'd128, 8'd128, 8'd128};
			{6'd0, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd23}: color = {8'd128, 8'd128, 8'd128};
			{6'd3, 6'd23}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd23}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd23}: color = {8'd64, 8'd64, 8'd64};
			{6'd6, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd23}: color = {8'd128, 8'd128, 8'd128};
			{6'd22, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd23}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd23}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd26, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd23}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd23}: color = {8'd192, 8'd192, 8'd128};
			{6'd46, 6'd23}: color = {8'd128, 8'd128, 8'd64};
			{6'd47, 6'd23}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd23}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd23}: color = {8'd64, 8'd64, 8'd0};
			{6'd50, 6'd23}: color = {8'd128, 8'd64, 8'd0};
			{6'd51, 6'd23}: color = {8'd128, 8'd128, 8'd64};
			{6'd52, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd23}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd23}: color = {8'd64, 8'd64, 8'd64};
			{6'd61, 6'd23}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd23}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd23}: color = {8'd128, 8'd128, 8'd128};
			{6'd0, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd24}: color = {8'd128, 8'd128, 8'd128};
			{6'd3, 6'd24}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd24}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd24}: color = {8'd192, 8'd128, 8'd128};
			{6'd22, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd24, 6'd24}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd24}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd24}: color = {8'd192, 8'd192, 8'd192};
			{6'd34, 6'd24}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd24}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd24}: color = {8'd192, 8'd128, 8'd128};
			{6'd46, 6'd24}: color = {8'd128, 8'd64, 8'd64};
			{6'd47, 6'd24}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd24}: color = {8'd64, 8'd64, 8'd0};
			{6'd49, 6'd24}: color = {8'd64, 8'd64, 8'd0};
			{6'd50, 6'd24}: color = {8'd128, 8'd64, 8'd64};
			{6'd51, 6'd24}: color = {8'd128, 8'd64, 8'd64};
			{6'd52, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd24}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd24}: color = {8'd128, 8'd128, 8'd128};
			{6'd62, 6'd24}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd24}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd25}: color = {8'd64, 8'd64, 8'd64};
			{6'd2, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd25}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd25}: color = {8'd64, 8'd64, 8'd64};
			{6'd20, 6'd25}: color = {8'd128, 8'd128, 8'd128};
			{6'd21, 6'd25}: color = {8'd64, 8'd64, 8'd0};
			{6'd22, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd25}: color = {8'd64, 8'd64, 8'd64};
			{6'd24, 6'd25}: color = {8'd128, 8'd128, 8'd128};
			{6'd25, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd34, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd25}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd25}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd25}: color = {8'd128, 8'd128, 8'd64};
			{6'd46, 6'd25}: color = {8'd128, 8'd64, 8'd0};
			{6'd47, 6'd25}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd25}: color = {8'd64, 8'd64, 8'd0};
			{6'd49, 6'd25}: color = {8'd128, 8'd64, 8'd0};
			{6'd50, 6'd25}: color = {8'd128, 8'd64, 8'd64};
			{6'd51, 6'd25}: color = {8'd128, 8'd64, 8'd0};
			{6'd52, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd25}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd25}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd25}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd26}: color = {8'd64, 8'd64, 8'd64};
			{6'd2, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd26}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd26}: color = {8'd192, 8'd128, 8'd128};
			{6'd21, 6'd26}: color = {8'd192, 8'd128, 8'd128};
			{6'd22, 6'd26}: color = {8'd192, 8'd128, 8'd64};
			{6'd23, 6'd26}: color = {8'd128, 8'd64, 8'd64};
			{6'd24, 6'd26}: color = {8'd128, 8'd64, 8'd0};
			{6'd25, 6'd26}: color = {8'd128, 8'd128, 8'd64};
			{6'd26, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd26}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd26}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd26}: color = {8'd128, 8'd64, 8'd0};
			{6'd46, 6'd26}: color = {8'd128, 8'd64, 8'd0};
			{6'd47, 6'd26}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd26}: color = {8'd64, 8'd64, 8'd0};
			{6'd49, 6'd26}: color = {8'd64, 8'd64, 8'd0};
			{6'd50, 6'd26}: color = {8'd128, 8'd128, 8'd64};
			{6'd51, 6'd26}: color = {8'd64, 8'd64, 8'd0};
			{6'd52, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd26}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd26}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd26}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd27}: color = {8'd64, 8'd64, 8'd64};
			{6'd2, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd27}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd21, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd22, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd27}: color = {8'd192, 8'd128, 8'd64};
			{6'd24, 6'd27}: color = {8'd192, 8'd64, 8'd64};
			{6'd25, 6'd27}: color = {8'd128, 8'd0, 8'd0};
			{6'd26, 6'd27}: color = {8'd128, 8'd128, 8'd64};
			{6'd27, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd27}: color = {8'd192, 8'd128, 8'd128};
			{6'd29, 6'd27}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd27}: color = {8'd192, 8'd128, 8'd128};
			{6'd31, 6'd27}: color = {8'd64, 8'd64, 8'd64};
			{6'd32, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd33, 6'd27}: color = {8'd64, 8'd64, 8'd0};
			{6'd34, 6'd27}: color = {8'd128, 8'd128, 8'd64};
			{6'd35, 6'd27}: color = {8'd192, 8'd128, 8'd128};
			{6'd36, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd39, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd27}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd27}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd27}: color = {8'd64, 8'd64, 8'd0};
			{6'd46, 6'd27}: color = {8'd128, 8'd64, 8'd0};
			{6'd47, 6'd27}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd27}: color = {8'd64, 8'd0, 8'd0};
			{6'd49, 6'd27}: color = {8'd64, 8'd64, 8'd0};
			{6'd50, 6'd27}: color = {8'd128, 8'd64, 8'd64};
			{6'd51, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd27}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd27}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd27}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd28}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd28}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd28}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd28}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd28}: color = {8'd128, 8'd128, 8'd128};
			{6'd20, 6'd28}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd28}: color = {8'd192, 8'd192, 8'd128};
			{6'd22, 6'd28}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd28}: color = {8'd192, 8'd128, 8'd128};
			{6'd24, 6'd28}: color = {8'd192, 8'd128, 8'd64};
			{6'd25, 6'd28}: color = {8'd128, 8'd64, 8'd0};
			{6'd26, 6'd28}: color = {8'd128, 8'd64, 8'd0};
			{6'd27, 6'd28}: color = {8'd192, 8'd128, 8'd64};
			{6'd28, 6'd28}: color = {8'd192, 8'd128, 8'd128};
			{6'd29, 6'd28}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd28}: color = {8'd128, 8'd64, 8'd64};
			{6'd31, 6'd28}: color = {8'd64, 8'd0, 8'd0};
			{6'd32, 6'd28}: color = {8'd128, 8'd64, 8'd0};
			{6'd33, 6'd28}: color = {8'd128, 8'd64, 8'd64};
			{6'd34, 6'd28}: color = {8'd128, 8'd64, 8'd64};
			{6'd35, 6'd28}: color = {8'd64, 8'd0, 8'd0};
			{6'd36, 6'd28}: color = {8'd192, 8'd128, 8'd128};
			{6'd37, 6'd28}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd28}: color = {8'd192, 8'd192, 8'd192};
			{6'd39, 6'd28}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd28}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd28}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd28}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd28}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd28}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd28}: color = {8'd64, 8'd64, 8'd0};
			{6'd46, 6'd28}: color = {8'd64, 8'd64, 8'd0};
			{6'd47, 6'd28}: color = {8'd64, 8'd64, 8'd0};
			{6'd48, 6'd28}: color = {8'd64, 8'd0, 8'd0};
			{6'd49, 6'd28}: color = {8'd128, 8'd64, 8'd64};
			{6'd50, 6'd28}: color = {8'd64, 8'd0, 8'd0};
			{6'd51, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd28}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd28}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd28}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd29}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd29}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd29}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd29}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd29}: color = {8'd192, 8'd192, 8'd128};
			{6'd21, 6'd29}: color = {8'd192, 8'd128, 8'd128};
			{6'd22, 6'd29}: color = {8'd192, 8'd128, 8'd128};
			{6'd23, 6'd29}: color = {8'd192, 8'd128, 8'd64};
			{6'd24, 6'd29}: color = {8'd128, 8'd64, 8'd64};
			{6'd25, 6'd29}: color = {8'd128, 8'd64, 8'd0};
			{6'd26, 6'd29}: color = {8'd128, 8'd64, 8'd0};
			{6'd27, 6'd29}: color = {8'd128, 8'd128, 8'd64};
			{6'd28, 6'd29}: color = {8'd192, 8'd128, 8'd128};
			{6'd29, 6'd29}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd29}: color = {8'd128, 8'd64, 8'd64};
			{6'd31, 6'd29}: color = {8'd128, 8'd64, 8'd0};
			{6'd32, 6'd29}: color = {8'd192, 8'd64, 8'd64};
			{6'd33, 6'd29}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd29}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd29}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd29}: color = {8'd128, 8'd64, 8'd64};
			{6'd37, 6'd29}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd29}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd29}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd29}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd29}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd29}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd29}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd29}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd29}: color = {8'd64, 8'd64, 8'd0};
			{6'd46, 6'd29}: color = {8'd64, 8'd64, 8'd0};
			{6'd47, 6'd29}: color = {8'd128, 8'd64, 8'd64};
			{6'd48, 6'd29}: color = {8'd128, 8'd64, 8'd64};
			{6'd49, 6'd29}: color = {8'd64, 8'd64, 8'd0};
			{6'd50, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd29}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd29}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd29}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd30}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd30}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd30}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd30}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd30}: color = {8'd128, 8'd128, 8'd128};
			{6'd21, 6'd30}: color = {8'd128, 8'd128, 8'd64};
			{6'd22, 6'd30}: color = {8'd64, 8'd64, 8'd64};
			{6'd23, 6'd30}: color = {8'd128, 8'd128, 8'd128};
			{6'd24, 6'd30}: color = {8'd128, 8'd128, 8'd128};
			{6'd25, 6'd30}: color = {8'd128, 8'd64, 8'd64};
			{6'd26, 6'd30}: color = {8'd128, 8'd64, 8'd0};
			{6'd27, 6'd30}: color = {8'd128, 8'd128, 8'd64};
			{6'd28, 6'd30}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd30}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd30}: color = {8'd192, 8'd64, 8'd64};
			{6'd31, 6'd30}: color = {8'd128, 8'd64, 8'd0};
			{6'd32, 6'd30}: color = {8'd128, 8'd64, 8'd0};
			{6'd33, 6'd30}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd30}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd30}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd30}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd30}: color = {8'd192, 8'd128, 8'd64};
			{6'd38, 6'd30}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd30}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd30}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd30}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd30}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd30}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd30}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd30}: color = {8'd128, 8'd64, 8'd64};
			{6'd46, 6'd30}: color = {8'd64, 8'd64, 8'd0};
			{6'd47, 6'd30}: color = {8'd128, 8'd128, 8'd64};
			{6'd48, 6'd30}: color = {8'd128, 8'd128, 8'd64};
			{6'd49, 6'd30}: color = {8'd128, 8'd128, 8'd128};
			{6'd50, 6'd30}: color = {8'd192, 8'd192, 8'd192};
			{6'd51, 6'd30}: color = {8'd64, 8'd64, 8'd64};
			{6'd52, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd30}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd30}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd30}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd31}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd31}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd31}: color = {8'd128, 8'd128, 8'd128};
			{6'd4, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd31}: color = {8'd64, 8'd0, 8'd0};
			{6'd19, 6'd31}: color = {8'd128, 8'd128, 8'd128};
			{6'd20, 6'd31}: color = {8'd128, 8'd128, 8'd128};
			{6'd21, 6'd31}: color = {8'd192, 8'd128, 8'd128};
			{6'd22, 6'd31}: color = {8'd192, 8'd128, 8'd128};
			{6'd23, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd24, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd31}: color = {8'd192, 8'd128, 8'd128};
			{6'd26, 6'd31}: color = {8'd192, 8'd128, 8'd64};
			{6'd27, 6'd31}: color = {8'd192, 8'd128, 8'd128};
			{6'd28, 6'd31}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd31}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd31}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd31}: color = {8'd128, 8'd64, 8'd64};
			{6'd32, 6'd31}: color = {8'd128, 8'd128, 8'd128};
			{6'd33, 6'd31}: color = {8'd64, 8'd64, 8'd64};
			{6'd34, 6'd31}: color = {8'd128, 8'd64, 8'd64};
			{6'd35, 6'd31}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd31}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd31}: color = {8'd192, 8'd128, 8'd64};
			{6'd38, 6'd31}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd44, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd45, 6'd31}: color = {8'd192, 8'd128, 8'd128};
			{6'd46, 6'd31}: color = {8'd64, 8'd0, 8'd0};
			{6'd47, 6'd31}: color = {8'd128, 8'd128, 8'd64};
			{6'd48, 6'd31}: color = {8'd192, 8'd192, 8'd128};
			{6'd49, 6'd31}: color = {8'd192, 8'd192, 8'd192};
			{6'd50, 6'd31}: color = {8'd192, 8'd192, 8'd192};
			{6'd51, 6'd31}: color = {8'd192, 8'd192, 8'd192};
			{6'd52, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd31}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd31}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd31}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd32}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd32}: color = {8'd128, 8'd128, 8'd128};
			{6'd4, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd32}: color = {8'd128, 8'd128, 8'd64};
			{6'd18, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd22, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd24, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd26, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd27, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd32, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd33, 6'd32}: color = {8'd128, 8'd128, 8'd64};
			{6'd34, 6'd32}: color = {8'd128, 8'd64, 8'd64};
			{6'd35, 6'd32}: color = {8'd64, 8'd64, 8'd64};
			{6'd36, 6'd32}: color = {8'd64, 8'd64, 8'd0};
			{6'd37, 6'd32}: color = {8'd128, 8'd128, 8'd64};
			{6'd38, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd32}: color = {8'd192, 8'd128, 8'd128};
			{6'd46, 6'd32}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd32}: color = {8'd192, 8'd128, 8'd64};
			{6'd48, 6'd32}: color = {8'd128, 8'd64, 8'd64};
			{6'd49, 6'd32}: color = {8'd64, 8'd0, 8'd0};
			{6'd50, 6'd32}: color = {8'd128, 8'd64, 8'd0};
			{6'd51, 6'd32}: color = {8'd192, 8'd192, 8'd128};
			{6'd52, 6'd32}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd32}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd32}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd32}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd33}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd33}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd33}: color = {8'd128, 8'd128, 8'd128};
			{6'd17, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd33}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd33}: color = {8'd192, 8'd128, 8'd128};
			{6'd26, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd33}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd33}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd33}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd33}: color = {8'd192, 8'd128, 8'd64};
			{6'd33, 6'd33}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd33}: color = {8'd192, 8'd64, 8'd0};
			{6'd35, 6'd33}: color = {8'd192, 8'd64, 8'd64};
			{6'd36, 6'd33}: color = {8'd128, 8'd64, 8'd64};
			{6'd37, 6'd33}: color = {8'd128, 8'd64, 8'd64};
			{6'd38, 6'd33}: color = {8'd192, 8'd128, 8'd64};
			{6'd39, 6'd33}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd33}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd33}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd33}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd33}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd33}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd33}: color = {8'd192, 8'd128, 8'd128};
			{6'd46, 6'd33}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd33}: color = {8'd128, 8'd64, 8'd64};
			{6'd48, 6'd33}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd33}: color = {8'd192, 8'd64, 8'd64};
			{6'd50, 6'd33}: color = {8'd128, 8'd64, 8'd0};
			{6'd51, 6'd33}: color = {8'd192, 8'd128, 8'd128};
			{6'd52, 6'd33}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd33}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd33}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd33}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd34}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd34}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd22, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd24, 6'd34}: color = {8'd192, 8'd128, 8'd128};
			{6'd25, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd34}: color = {8'd192, 8'd128, 8'd128};
			{6'd35, 6'd34}: color = {8'd192, 8'd128, 8'd128};
			{6'd36, 6'd34}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd34}: color = {8'd192, 8'd128, 8'd64};
			{6'd38, 6'd34}: color = {8'd192, 8'd128, 8'd64};
			{6'd39, 6'd34}: color = {8'd192, 8'd128, 8'd64};
			{6'd40, 6'd34}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd34}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd34}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd34}: color = {8'd192, 8'd128, 8'd128};
			{6'd46, 6'd34}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd34}: color = {8'd64, 8'd0, 8'd0};
			{6'd48, 6'd34}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd34}: color = {8'd192, 8'd128, 8'd64};
			{6'd50, 6'd34}: color = {8'd128, 8'd64, 8'd0};
			{6'd51, 6'd34}: color = {8'd192, 8'd192, 8'd128};
			{6'd52, 6'd34}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd34}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd34}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd34}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd35}: color = {8'd128, 8'd128, 8'd128};
			{6'd2, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd35}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd17, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd21, 6'd35}: color = {8'd192, 8'd128, 8'd64};
			{6'd22, 6'd35}: color = {8'd128, 8'd64, 8'd64};
			{6'd23, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd24, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd31, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd32, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd33, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd35}: color = {8'd192, 8'd128, 8'd64};
			{6'd39, 6'd35}: color = {8'd192, 8'd128, 8'd64};
			{6'd40, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd35}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd35}: color = {8'd192, 8'd128, 8'd128};
			{6'd46, 6'd35}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd35}: color = {8'd128, 8'd0, 8'd0};
			{6'd48, 6'd35}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd35}: color = {8'd128, 8'd64, 8'd64};
			{6'd50, 6'd35}: color = {8'd192, 8'd128, 8'd64};
			{6'd51, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd52, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd35}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd35}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd35}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd36}: color = {8'd64, 8'd64, 8'd64};
			{6'd2, 6'd36}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd36}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd36}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd36}: color = {8'd128, 8'd128, 8'd128};
			{6'd17, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd18, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd19, 6'd36}: color = {8'd192, 8'd128, 8'd64};
			{6'd20, 6'd36}: color = {8'd192, 8'd64, 8'd64};
			{6'd21, 6'd36}: color = {8'd128, 8'd64, 8'd0};
			{6'd22, 6'd36}: color = {8'd128, 8'd64, 8'd64};
			{6'd23, 6'd36}: color = {8'd128, 8'd128, 8'd64};
			{6'd24, 6'd36}: color = {8'd192, 8'd128, 8'd64};
			{6'd25, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd26, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd31, 6'd36}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd36}: color = {8'd128, 8'd64, 8'd64};
			{6'd33, 6'd36}: color = {8'd192, 8'd64, 8'd64};
			{6'd34, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd36}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd36}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd36}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd36}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd36}: color = {8'd192, 8'd128, 8'd64};
			{6'd46, 6'd36}: color = {8'd128, 8'd64, 8'd64};
			{6'd47, 6'd36}: color = {8'd128, 8'd0, 8'd0};
			{6'd48, 6'd36}: color = {8'd128, 8'd64, 8'd0};
			{6'd49, 6'd36}: color = {8'd128, 8'd64, 8'd64};
			{6'd50, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd51, 6'd36}: color = {8'd192, 8'd128, 8'd128};
			{6'd52, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd36}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd36}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd36}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd36}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd37}: color = {8'd64, 8'd64, 8'd64};
			{6'd2, 6'd37}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd37}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd37}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd37}: color = {8'd128, 8'd128, 8'd64};
			{6'd17, 6'd37}: color = {8'd192, 8'd192, 8'd128};
			{6'd18, 6'd37}: color = {8'd192, 8'd128, 8'd64};
			{6'd19, 6'd37}: color = {8'd192, 8'd64, 8'd64};
			{6'd20, 6'd37}: color = {8'd128, 8'd64, 8'd0};
			{6'd21, 6'd37}: color = {8'd128, 8'd64, 8'd64};
			{6'd22, 6'd37}: color = {8'd192, 8'd128, 8'd128};
			{6'd23, 6'd37}: color = {8'd192, 8'd128, 8'd64};
			{6'd24, 6'd37}: color = {8'd128, 8'd64, 8'd0};
			{6'd25, 6'd37}: color = {8'd128, 8'd64, 8'd0};
			{6'd26, 6'd37}: color = {8'd192, 8'd64, 8'd64};
			{6'd27, 6'd37}: color = {8'd64, 8'd64, 8'd64};
			{6'd28, 6'd37}: color = {8'd64, 8'd64, 8'd0};
			{6'd29, 6'd37}: color = {8'd128, 8'd64, 8'd64};
			{6'd30, 6'd37}: color = {8'd128, 8'd64, 8'd64};
			{6'd31, 6'd37}: color = {8'd128, 8'd64, 8'd64};
			{6'd32, 6'd37}: color = {8'd128, 8'd128, 8'd64};
			{6'd33, 6'd37}: color = {8'd192, 8'd64, 8'd64};
			{6'd34, 6'd37}: color = {8'd128, 8'd64, 8'd64};
			{6'd35, 6'd37}: color = {8'd192, 8'd128, 8'd128};
			{6'd36, 6'd37}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd37}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd37}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd37}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd37}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd37}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd37}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd37}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd37}: color = {8'd192, 8'd128, 8'd128};
			{6'd45, 6'd37}: color = {8'd192, 8'd128, 8'd64};
			{6'd46, 6'd37}: color = {8'd128, 8'd0, 8'd0};
			{6'd47, 6'd37}: color = {8'd128, 8'd0, 8'd0};
			{6'd48, 6'd37}: color = {8'd128, 8'd64, 8'd64};
			{6'd49, 6'd37}: color = {8'd128, 8'd128, 8'd64};
			{6'd50, 6'd37}: color = {8'd192, 8'd192, 8'd128};
			{6'd51, 6'd37}: color = {8'd64, 8'd64, 8'd64};
			{6'd52, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd37}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd37}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd37}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd37}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd38}: color = {8'd64, 8'd64, 8'd64};
			{6'd2, 6'd38}: color = {8'd192, 8'd192, 8'd192};
			{6'd3, 6'd38}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd38}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd38}: color = {8'd64, 8'd64, 8'd64};
			{6'd17, 6'd38}: color = {8'd192, 8'd192, 8'd128};
			{6'd18, 6'd38}: color = {8'd192, 8'd64, 8'd64};
			{6'd19, 6'd38}: color = {8'd128, 8'd64, 8'd0};
			{6'd20, 6'd38}: color = {8'd128, 8'd64, 8'd64};
			{6'd21, 6'd38}: color = {8'd192, 8'd128, 8'd128};
			{6'd22, 6'd38}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd38}: color = {8'd192, 8'd192, 8'd128};
			{6'd24, 6'd38}: color = {8'd192, 8'd64, 8'd64};
			{6'd25, 6'd38}: color = {8'd128, 8'd64, 8'd0};
			{6'd26, 6'd38}: color = {8'd64, 8'd0, 8'd0};
			{6'd27, 6'd38}: color = {8'd64, 8'd0, 8'd0};
			{6'd28, 6'd38}: color = {8'd64, 8'd0, 8'd0};
			{6'd29, 6'd38}: color = {8'd128, 8'd0, 8'd0};
			{6'd30, 6'd38}: color = {8'd128, 8'd0, 8'd0};
			{6'd31, 6'd38}: color = {8'd128, 8'd64, 8'd64};
			{6'd32, 6'd38}: color = {8'd192, 8'd128, 8'd128};
			{6'd33, 6'd38}: color = {8'd192, 8'd128, 8'd128};
			{6'd34, 6'd38}: color = {8'd128, 8'd64, 8'd0};
			{6'd35, 6'd38}: color = {8'd128, 8'd64, 8'd0};
			{6'd36, 6'd38}: color = {8'd192, 8'd64, 8'd64};
			{6'd37, 6'd38}: color = {8'd192, 8'd128, 8'd64};
			{6'd38, 6'd38}: color = {8'd192, 8'd128, 8'd64};
			{6'd39, 6'd38}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd38}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd38}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd38}: color = {8'd192, 8'd192, 8'd128};
			{6'd43, 6'd38}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd38}: color = {8'd192, 8'd128, 8'd64};
			{6'd45, 6'd38}: color = {8'd192, 8'd128, 8'd64};
			{6'd46, 6'd38}: color = {8'd128, 8'd64, 8'd64};
			{6'd47, 6'd38}: color = {8'd128, 8'd64, 8'd64};
			{6'd48, 6'd38}: color = {8'd192, 8'd128, 8'd64};
			{6'd49, 6'd38}: color = {8'd192, 8'd128, 8'd64};
			{6'd50, 6'd38}: color = {8'd192, 8'd128, 8'd128};
			{6'd51, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd38}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd38}: color = {8'd128, 8'd128, 8'd128};
			{6'd62, 6'd38}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd38}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd39}: color = {8'd128, 8'd128, 8'd128};
			{6'd3, 6'd39}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd39}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd39}: color = {8'd128, 8'd128, 8'd128};
			{6'd17, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd18, 6'd39}: color = {8'd128, 8'd64, 8'd64};
			{6'd19, 6'd39}: color = {8'd128, 8'd64, 8'd64};
			{6'd20, 6'd39}: color = {8'd192, 8'd128, 8'd128};
			{6'd21, 6'd39}: color = {8'd192, 8'd128, 8'd128};
			{6'd22, 6'd39}: color = {8'd192, 8'd128, 8'd128};
			{6'd23, 6'd39}: color = {8'd192, 8'd128, 8'd128};
			{6'd24, 6'd39}: color = {8'd192, 8'd128, 8'd64};
			{6'd25, 6'd39}: color = {8'd192, 8'd64, 8'd0};
			{6'd26, 6'd39}: color = {8'd192, 8'd64, 8'd0};
			{6'd27, 6'd39}: color = {8'd192, 8'd64, 8'd0};
			{6'd28, 6'd39}: color = {8'd128, 8'd64, 8'd0};
			{6'd29, 6'd39}: color = {8'd128, 8'd64, 8'd0};
			{6'd30, 6'd39}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd39}: color = {8'd192, 8'd64, 8'd64};
			{6'd36, 6'd39}: color = {8'd128, 8'd64, 8'd0};
			{6'd37, 6'd39}: color = {8'd128, 8'd64, 8'd0};
			{6'd38, 6'd39}: color = {8'd192, 8'd64, 8'd64};
			{6'd39, 6'd39}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd39}: color = {8'd192, 8'd128, 8'd128};
			{6'd43, 6'd39}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd39}: color = {8'd192, 8'd128, 8'd64};
			{6'd45, 6'd39}: color = {8'd192, 8'd128, 8'd64};
			{6'd46, 6'd39}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd39}: color = {8'd192, 8'd128, 8'd64};
			{6'd48, 6'd39}: color = {8'd128, 8'd128, 8'd64};
			{6'd49, 6'd39}: color = {8'd192, 8'd192, 8'd128};
			{6'd50, 6'd39}: color = {8'd64, 8'd64, 8'd64};
			{6'd51, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd39}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd39}: color = {8'd128, 8'd128, 8'd128};
			{6'd62, 6'd39}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd39}: color = {8'd192, 8'd192, 8'd192};
			{6'd0, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd40}: color = {8'd128, 8'd128, 8'd128};
			{6'd3, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd40}: color = {8'd64, 8'd64, 8'd64};
			{6'd6, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd40}: color = {8'd128, 8'd128, 8'd128};
			{6'd17, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd40}: color = {8'd192, 8'd192, 8'd128};
			{6'd19, 6'd40}: color = {8'd192, 8'd128, 8'd128};
			{6'd20, 6'd40}: color = {8'd64, 8'd64, 8'd64};
			{6'd21, 6'd40}: color = {8'd64, 8'd64, 8'd64};
			{6'd22, 6'd40}: color = {8'd128, 8'd64, 8'd64};
			{6'd23, 6'd40}: color = {8'd128, 8'd64, 8'd64};
			{6'd24, 6'd40}: color = {8'd128, 8'd64, 8'd64};
			{6'd25, 6'd40}: color = {8'd128, 8'd0, 8'd0};
			{6'd26, 6'd40}: color = {8'd128, 8'd0, 8'd0};
			{6'd27, 6'd40}: color = {8'd128, 8'd0, 8'd0};
			{6'd28, 6'd40}: color = {8'd192, 8'd64, 8'd0};
			{6'd29, 6'd40}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd32, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd33, 6'd40}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd40}: color = {8'd128, 8'd64, 8'd64};
			{6'd35, 6'd40}: color = {8'd128, 8'd64, 8'd64};
			{6'd36, 6'd40}: color = {8'd192, 8'd128, 8'd128};
			{6'd37, 6'd40}: color = {8'd128, 8'd64, 8'd64};
			{6'd38, 6'd40}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd40}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd40}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd40}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd40}: color = {8'd192, 8'd128, 8'd128};
			{6'd43, 6'd40}: color = {8'd192, 8'd128, 8'd128};
			{6'd44, 6'd40}: color = {8'd192, 8'd128, 8'd64};
			{6'd45, 6'd40}: color = {8'd192, 8'd64, 8'd64};
			{6'd46, 6'd40}: color = {8'd192, 8'd128, 8'd64};
			{6'd47, 6'd40}: color = {8'd192, 8'd128, 8'd64};
			{6'd48, 6'd40}: color = {8'd192, 8'd192, 8'd128};
			{6'd49, 6'd40}: color = {8'd64, 8'd64, 8'd64};
			{6'd50, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd40}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd40}: color = {8'd64, 8'd64, 8'd64};
			{6'd61, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd40}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd40}: color = {8'd128, 8'd128, 8'd128};
			{6'd0, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd41}: color = {8'd64, 8'd64, 8'd64};
			{6'd3, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd4, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd41}: color = {8'd128, 8'd128, 8'd128};
			{6'd6, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd21, 6'd41}: color = {8'd128, 8'd128, 8'd128};
			{6'd22, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd26, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd27, 6'd41}: color = {8'd128, 8'd64, 8'd64};
			{6'd28, 6'd41}: color = {8'd128, 8'd64, 8'd0};
			{6'd29, 6'd41}: color = {8'd192, 8'd64, 8'd64};
			{6'd30, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd31, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd32, 6'd41}: color = {8'd128, 8'd128, 8'd128};
			{6'd33, 6'd41}: color = {8'd64, 8'd64, 8'd64};
			{6'd34, 6'd41}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd36, 6'd41}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd41}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd41}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd41}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd41}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd41}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd43, 6'd41}: color = {8'd192, 8'd128, 8'd64};
			{6'd44, 6'd41}: color = {8'd64, 8'd64, 8'd0};
			{6'd45, 6'd41}: color = {8'd192, 8'd128, 8'd64};
			{6'd46, 6'd41}: color = {8'd192, 8'd192, 8'd128};
			{6'd47, 6'd41}: color = {8'd192, 8'd128, 8'd128};
			{6'd48, 6'd41}: color = {8'd64, 8'd64, 8'd64};
			{6'd49, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd41}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd41}: color = {8'd64, 8'd64, 8'd64};
			{6'd61, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd41}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd41}: color = {8'd64, 8'd64, 8'd64};
			{6'd0, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd42}: color = {8'd128, 8'd128, 8'd128};
			{6'd4, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd42}: color = {8'd128, 8'd128, 8'd128};
			{6'd6, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd19, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd20, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd21, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd42}: color = {8'd128, 8'd128, 8'd128};
			{6'd30, 6'd42}: color = {8'd128, 8'd64, 8'd64};
			{6'd31, 6'd42}: color = {8'd64, 8'd0, 8'd0};
			{6'd32, 6'd42}: color = {8'd128, 8'd64, 8'd64};
			{6'd33, 6'd42}: color = {8'd192, 8'd128, 8'd128};
			{6'd34, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd42}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd42}: color = {8'd192, 8'd128, 8'd128};
			{6'd43, 6'd42}: color = {8'd128, 8'd64, 8'd0};
			{6'd44, 6'd42}: color = {8'd64, 8'd64, 8'd0};
			{6'd45, 6'd42}: color = {8'd64, 8'd64, 8'd64};
			{6'd46, 6'd42}: color = {8'd64, 8'd64, 8'd64};
			{6'd47, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd42}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd42}: color = {8'd128, 8'd128, 8'd128};
			{6'd61, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd42}: color = {8'd192, 8'd192, 8'd192};
			{6'd63, 6'd42}: color = {8'd64, 8'd64, 8'd64};
			{6'd0, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd43}: color = {8'd128, 8'd128, 8'd128};
			{6'd4, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd43}: color = {8'd64, 8'd64, 8'd64};
			{6'd7, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd43}: color = {8'd128, 8'd128, 8'd128};
			{6'd17, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd43}: color = {8'd192, 8'd128, 8'd128};
			{6'd19, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd20, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd21, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd22, 6'd43}: color = {8'd192, 8'd128, 8'd128};
			{6'd23, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd43}: color = {8'd128, 8'd128, 8'd128};
			{6'd31, 6'd43}: color = {8'd192, 8'd128, 8'd128};
			{6'd32, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd43}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd43}: color = {8'd192, 8'd128, 8'd64};
			{6'd43, 6'd43}: color = {8'd64, 8'd64, 8'd0};
			{6'd44, 6'd43}: color = {8'd64, 8'd64, 8'd64};
			{6'd45, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd43}: color = {8'd64, 8'd64, 8'd64};
			{6'd60, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd43}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd43}: color = {8'd128, 8'd128, 8'd128};
			{6'd63, 6'd43}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd44}: color = {8'd64, 8'd64, 8'd64};
			{6'd4, 6'd44}: color = {8'd192, 8'd192, 8'd192};
			{6'd5, 6'd44}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd44}: color = {8'd128, 8'd128, 8'd128};
			{6'd7, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd44}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd19, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd20, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd21, 6'd44}: color = {8'd192, 8'd128, 8'd64};
			{6'd22, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd23, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd24, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd25, 6'd44}: color = {8'd192, 8'd128, 8'd64};
			{6'd26, 6'd44}: color = {8'd192, 8'd128, 8'd64};
			{6'd27, 6'd44}: color = {8'd192, 8'd64, 8'd64};
			{6'd28, 6'd44}: color = {8'd192, 8'd128, 8'd64};
			{6'd29, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd31, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd44}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd44}: color = {8'd192, 8'd128, 8'd128};
			{6'd42, 6'd44}: color = {8'd128, 8'd64, 8'd64};
			{6'd43, 6'd44}: color = {8'd64, 8'd64, 8'd0};
			{6'd44, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd44}: color = {8'd128, 8'd128, 8'd128};
			{6'd60, 6'd44}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd44}: color = {8'd192, 8'd192, 8'd192};
			{6'd62, 6'd44}: color = {8'd64, 8'd64, 8'd64};
			{6'd63, 6'd44}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd45}: color = {8'd128, 8'd128, 8'd128};
			{6'd5, 6'd45}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd45}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd45}: color = {8'd64, 8'd64, 8'd64};
			{6'd8, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd45}: color = {8'd128, 8'd128, 8'd128};
			{6'd18, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd19, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd20, 6'd45}: color = {8'd192, 8'd128, 8'd128};
			{6'd21, 6'd45}: color = {8'd192, 8'd128, 8'd64};
			{6'd22, 6'd45}: color = {8'd128, 8'd128, 8'd64};
			{6'd23, 6'd45}: color = {8'd192, 8'd128, 8'd128};
			{6'd24, 6'd45}: color = {8'd192, 8'd128, 8'd128};
			{6'd25, 6'd45}: color = {8'd192, 8'd128, 8'd64};
			{6'd26, 6'd45}: color = {8'd192, 8'd64, 8'd0};
			{6'd27, 6'd45}: color = {8'd192, 8'd64, 8'd0};
			{6'd28, 6'd45}: color = {8'd128, 8'd64, 8'd64};
			{6'd29, 6'd45}: color = {8'd192, 8'd128, 8'd128};
			{6'd30, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd45}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd45}: color = {8'd192, 8'd128, 8'd128};
			{6'd42, 6'd45}: color = {8'd128, 8'd128, 8'd64};
			{6'd43, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd45}: color = {8'd64, 8'd64, 8'd64};
			{6'd59, 6'd45}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd45}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd45}: color = {8'd128, 8'd128, 8'd128};
			{6'd62, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd45}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd46}: color = {8'd64, 8'd64, 8'd64};
			{6'd5, 6'd46}: color = {8'd192, 8'd192, 8'd192};
			{6'd6, 6'd46}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd46}: color = {8'd128, 8'd128, 8'd128};
			{6'd8, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd46}: color = {8'd192, 8'd128, 8'd128};
			{6'd19, 6'd46}: color = {8'd192, 8'd128, 8'd128};
			{6'd20, 6'd46}: color = {8'd192, 8'd128, 8'd64};
			{6'd21, 6'd46}: color = {8'd192, 8'd128, 8'd64};
			{6'd22, 6'd46}: color = {8'd192, 8'd128, 8'd64};
			{6'd23, 6'd46}: color = {8'd128, 8'd64, 8'd64};
			{6'd24, 6'd46}: color = {8'd128, 8'd64, 8'd64};
			{6'd25, 6'd46}: color = {8'd128, 8'd64, 8'd64};
			{6'd26, 6'd46}: color = {8'd128, 8'd64, 8'd64};
			{6'd27, 6'd46}: color = {8'd128, 8'd128, 8'd128};
			{6'd28, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd46}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd46}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd46}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd46}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd46}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd46}: color = {8'd64, 8'd64, 8'd64};
			{6'd43, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd46}: color = {8'd128, 8'd128, 8'd128};
			{6'd59, 6'd46}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd46}: color = {8'd192, 8'd192, 8'd192};
			{6'd61, 6'd46}: color = {8'd64, 8'd64, 8'd64};
			{6'd62, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd46}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd47}: color = {8'd128, 8'd128, 8'd128};
			{6'd6, 6'd47}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd47}: color = {8'd192, 8'd192, 8'd192};
			{6'd8, 6'd47}: color = {8'd128, 8'd128, 8'd128};
			{6'd9, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd47}: color = {8'd64, 8'd64, 8'd64};
			{6'd17, 6'd47}: color = {8'd192, 8'd128, 8'd128};
			{6'd18, 6'd47}: color = {8'd192, 8'd128, 8'd128};
			{6'd19, 6'd47}: color = {8'd192, 8'd128, 8'd128};
			{6'd20, 6'd47}: color = {8'd192, 8'd128, 8'd128};
			{6'd21, 6'd47}: color = {8'd192, 8'd128, 8'd64};
			{6'd22, 6'd47}: color = {8'd192, 8'd128, 8'd64};
			{6'd23, 6'd47}: color = {8'd192, 8'd128, 8'd64};
			{6'd24, 6'd47}: color = {8'd192, 8'd128, 8'd64};
			{6'd25, 6'd47}: color = {8'd192, 8'd128, 8'd64};
			{6'd26, 6'd47}: color = {8'd192, 8'd128, 8'd64};
			{6'd27, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd47}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd38, 6'd47}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd47}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd47}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd47}: color = {8'd128, 8'd128, 8'd128};
			{6'd42, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd47}: color = {8'd64, 8'd64, 8'd64};
			{6'd58, 6'd47}: color = {8'd192, 8'd192, 8'd192};
			{6'd59, 6'd47}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd47}: color = {8'd128, 8'd128, 8'd128};
			{6'd61, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd47}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd48}: color = {8'd64, 8'd64, 8'd64};
			{6'd6, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd7, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd8, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd48}: color = {8'd64, 8'd64, 8'd64};
			{6'd10, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd48}: color = {8'd64, 8'd64, 8'd64};
			{6'd16, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd18, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd19, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd20, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd23, 6'd48}: color = {8'd192, 8'd128, 8'd128};
			{6'd24, 6'd48}: color = {8'd192, 8'd128, 8'd128};
			{6'd25, 6'd48}: color = {8'd192, 8'd128, 8'd128};
			{6'd26, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd35, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd36, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd48}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd48}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd48}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd48}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd48}: color = {8'd64, 8'd64, 8'd64};
			{6'd42, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd48}: color = {8'd64, 8'd64, 8'd64};
			{6'd57, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd58, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd59, 6'd48}: color = {8'd192, 8'd192, 8'd192};
			{6'd60, 6'd48}: color = {8'd64, 8'd64, 8'd64};
			{6'd61, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd48}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd49}: color = {8'd64, 8'd64, 8'd64};
			{6'd7, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd8, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd49}: color = {8'd128, 8'd128, 8'd128};
			{6'd10, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd49}: color = {8'd128, 8'd128, 8'd128};
			{6'd16, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd17, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd18, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd26, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd32, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd34, 6'd49}: color = {8'd192, 8'd128, 8'd128};
			{6'd35, 6'd49}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd49}: color = {8'd192, 8'd128, 8'd128};
			{6'd37, 6'd49}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd49}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd49}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd49}: color = {8'd64, 8'd0, 8'd0};
			{6'd42, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd49}: color = {8'd128, 8'd128, 8'd128};
			{6'd57, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd58, 6'd49}: color = {8'd192, 8'd192, 8'd192};
			{6'd59, 6'd49}: color = {8'd128, 8'd128, 8'd128};
			{6'd60, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd49}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd50}: color = {8'd128, 8'd128, 8'd128};
			{6'd8, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd10, 6'd50}: color = {8'd128, 8'd128, 8'd128};
			{6'd11, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd16, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd17, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd18, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd27, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd29, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd30, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd31, 6'd50}: color = {8'd192, 8'd128, 8'd128};
			{6'd32, 6'd50}: color = {8'd192, 8'd128, 8'd64};
			{6'd33, 6'd50}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd50}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd50}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd50}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd50}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd50}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd50}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd50}: color = {8'd128, 8'd128, 8'd128};
			{6'd56, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd57, 6'd50}: color = {8'd192, 8'd192, 8'd192};
			{6'd58, 6'd50}: color = {8'd128, 8'd128, 8'd128};
			{6'd59, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd50}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd51}: color = {8'd64, 8'd64, 8'd64};
			{6'd8, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd9, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd10, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd11, 6'd51}: color = {8'd128, 8'd128, 8'd128};
			{6'd12, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd16, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd17, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd18, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd19, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd20, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd21, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd24, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd25, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd26, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd27, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd28, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd29, 6'd51}: color = {8'd192, 8'd128, 8'd64};
			{6'd30, 6'd51}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd51}: color = {8'd192, 8'd64, 8'd0};
			{6'd32, 6'd51}: color = {8'd192, 8'd64, 8'd0};
			{6'd33, 6'd51}: color = {8'd192, 8'd64, 8'd64};
			{6'd34, 6'd51}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd51}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd51}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd51}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd51}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd51}: color = {8'd64, 8'd64, 8'd64};
			{6'd55, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd56, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd57, 6'd51}: color = {8'd192, 8'd192, 8'd192};
			{6'd58, 6'd51}: color = {8'd64, 8'd64, 8'd64};
			{6'd59, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd51}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd52}: color = {8'd64, 8'd64, 8'd64};
			{6'd9, 6'd52}: color = {8'd192, 8'd192, 8'd192};
			{6'd10, 6'd52}: color = {8'd192, 8'd192, 8'd192};
			{6'd11, 6'd52}: color = {8'd192, 8'd192, 8'd192};
			{6'd12, 6'd52}: color = {8'd128, 8'd128, 8'd128};
			{6'd13, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd52}: color = {8'd192, 8'd128, 8'd128};
			{6'd17, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd18, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd19, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd20, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd21, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd22, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd23, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd24, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd25, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd26, 6'd52}: color = {8'd128, 8'd128, 8'd64};
			{6'd27, 6'd52}: color = {8'd192, 8'd64, 8'd64};
			{6'd28, 6'd52}: color = {8'd192, 8'd64, 8'd64};
			{6'd29, 6'd52}: color = {8'd192, 8'd64, 8'd0};
			{6'd30, 6'd52}: color = {8'd192, 8'd64, 8'd0};
			{6'd31, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd33, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd52}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd52}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd52}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd52}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd52}: color = {8'd192, 8'd128, 8'd128};
			{6'd41, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd52}: color = {8'd64, 8'd64, 8'd64};
			{6'd54, 6'd52}: color = {8'd192, 8'd192, 8'd192};
			{6'd55, 6'd52}: color = {8'd192, 8'd192, 8'd192};
			{6'd56, 6'd52}: color = {8'd192, 8'd192, 8'd192};
			{6'd57, 6'd52}: color = {8'd64, 8'd64, 8'd64};
			{6'd58, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd52}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd53}: color = {8'd64, 8'd64, 8'd64};
			{6'd10, 6'd53}: color = {8'd192, 8'd192, 8'd192};
			{6'd11, 6'd53}: color = {8'd192, 8'd192, 8'd192};
			{6'd12, 6'd53}: color = {8'd192, 8'd192, 8'd192};
			{6'd13, 6'd53}: color = {8'd128, 8'd128, 8'd128};
			{6'd14, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd53}: color = {8'd128, 8'd64, 8'd64};
			{6'd18, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd19, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd20, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd21, 6'd53}: color = {8'd192, 8'd64, 8'd64};
			{6'd22, 6'd53}: color = {8'd192, 8'd64, 8'd0};
			{6'd23, 6'd53}: color = {8'd128, 8'd64, 8'd0};
			{6'd24, 6'd53}: color = {8'd128, 8'd64, 8'd0};
			{6'd25, 6'd53}: color = {8'd128, 8'd64, 8'd64};
			{6'd26, 6'd53}: color = {8'd192, 8'd64, 8'd64};
			{6'd27, 6'd53}: color = {8'd192, 8'd64, 8'd64};
			{6'd28, 6'd53}: color = {8'd192, 8'd64, 8'd64};
			{6'd29, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd30, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd33, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd53}: color = {8'd192, 8'd128, 8'd64};
			{6'd37, 6'd53}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd53}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd53}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd53}: color = {8'd128, 8'd128, 8'd64};
			{6'd41, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd53}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd53}: color = {8'd192, 8'd192, 8'd192};
			{6'd54, 6'd53}: color = {8'd192, 8'd192, 8'd192};
			{6'd55, 6'd53}: color = {8'd192, 8'd192, 8'd192};
			{6'd56, 6'd53}: color = {8'd64, 8'd64, 8'd64};
			{6'd57, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd53}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd54}: color = {8'd64, 8'd64, 8'd64};
			{6'd11, 6'd54}: color = {8'd192, 8'd192, 8'd192};
			{6'd12, 6'd54}: color = {8'd192, 8'd192, 8'd192};
			{6'd13, 6'd54}: color = {8'd192, 8'd192, 8'd192};
			{6'd14, 6'd54}: color = {8'd128, 8'd128, 8'd128};
			{6'd15, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd54}: color = {8'd64, 8'd0, 8'd0};
			{6'd20, 6'd54}: color = {8'd64, 8'd64, 8'd0};
			{6'd21, 6'd54}: color = {8'd128, 8'd64, 8'd64};
			{6'd22, 6'd54}: color = {8'd128, 8'd64, 8'd64};
			{6'd23, 6'd54}: color = {8'd128, 8'd64, 8'd64};
			{6'd24, 6'd54}: color = {8'd192, 8'd64, 8'd64};
			{6'd25, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd26, 6'd54}: color = {8'd192, 8'd64, 8'd64};
			{6'd27, 6'd54}: color = {8'd192, 8'd64, 8'd64};
			{6'd28, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd29, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd30, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd33, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd54}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd54}: color = {8'd192, 8'd128, 8'd128};
			{6'd37, 6'd54}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd54}: color = {8'd192, 8'd128, 8'd128};
			{6'd39, 6'd54}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd54}: color = {8'd128, 8'd128, 8'd128};
			{6'd52, 6'd54}: color = {8'd192, 8'd192, 8'd192};
			{6'd53, 6'd54}: color = {8'd192, 8'd192, 8'd192};
			{6'd54, 6'd54}: color = {8'd192, 8'd192, 8'd192};
			{6'd55, 6'd54}: color = {8'd128, 8'd128, 8'd128};
			{6'd56, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd54}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd55}: color = {8'd64, 8'd64, 8'd64};
			{6'd12, 6'd55}: color = {8'd192, 8'd192, 8'd192};
			{6'd13, 6'd55}: color = {8'd192, 8'd192, 8'd192};
			{6'd14, 6'd55}: color = {8'd192, 8'd192, 8'd192};
			{6'd15, 6'd55}: color = {8'd128, 8'd128, 8'd128};
			{6'd16, 6'd55}: color = {8'd64, 8'd64, 8'd64};
			{6'd17, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd55}: color = {8'd128, 8'd128, 8'd128};
			{6'd24, 6'd55}: color = {8'd192, 8'd128, 8'd128};
			{6'd25, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd26, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd27, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd28, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd29, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd30, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd33, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd34, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd55}: color = {8'd192, 8'd128, 8'd64};
			{6'd36, 6'd55}: color = {8'd192, 8'd128, 8'd128};
			{6'd37, 6'd55}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd55}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd55}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd55}: color = {8'd64, 8'd64, 8'd64};
			{6'd41, 6'd55}: color = {8'd64, 8'd64, 8'd64};
			{6'd42, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd55}: color = {8'd64, 8'd64, 8'd64};
			{6'd50, 6'd55}: color = {8'd128, 8'd128, 8'd128};
			{6'd51, 6'd55}: color = {8'd192, 8'd192, 8'd192};
			{6'd52, 6'd55}: color = {8'd192, 8'd192, 8'd192};
			{6'd53, 6'd55}: color = {8'd192, 8'd192, 8'd192};
			{6'd54, 6'd55}: color = {8'd64, 8'd64, 8'd64};
			{6'd55, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd55}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd56}: color = {8'd64, 8'd64, 8'd64};
			{6'd13, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd14, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd15, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd16, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd56}: color = {8'd128, 8'd128, 8'd128};
			{6'd18, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd56}: color = {8'd64, 8'd64, 8'd64};
			{6'd25, 6'd56}: color = {8'd128, 8'd128, 8'd128};
			{6'd26, 6'd56}: color = {8'd192, 8'd128, 8'd128};
			{6'd27, 6'd56}: color = {8'd192, 8'd128, 8'd64};
			{6'd28, 6'd56}: color = {8'd192, 8'd128, 8'd64};
			{6'd29, 6'd56}: color = {8'd192, 8'd128, 8'd64};
			{6'd30, 6'd56}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd56}: color = {8'd192, 8'd128, 8'd64};
			{6'd32, 6'd56}: color = {8'd192, 8'd128, 8'd128};
			{6'd33, 6'd56}: color = {8'd192, 8'd128, 8'd128};
			{6'd34, 6'd56}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd56}: color = {8'd192, 8'd128, 8'd128};
			{6'd36, 6'd56}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd56}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd56}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd56}: color = {8'd192, 8'd128, 8'd128};
			{6'd40, 6'd56}: color = {8'd192, 8'd192, 8'd128};
			{6'd41, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd42, 6'd56}: color = {8'd0, 8'd0, 8'd64};
			{6'd43, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd56}: color = {8'd64, 8'd64, 8'd64};
			{6'd49, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd50, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd51, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd52, 6'd56}: color = {8'd192, 8'd192, 8'd192};
			{6'd53, 6'd56}: color = {8'd64, 8'd64, 8'd64};
			{6'd54, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd56}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd57}: color = {8'd64, 8'd64, 8'd64};
			{6'd14, 6'd57}: color = {8'd128, 8'd128, 8'd128};
			{6'd15, 6'd57}: color = {8'd192, 8'd192, 8'd192};
			{6'd16, 6'd57}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd57}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd57}: color = {8'd128, 8'd128, 8'd128};
			{6'd19, 6'd57}: color = {8'd64, 8'd64, 8'd64};
			{6'd20, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd57}: color = {8'd64, 8'd64, 8'd64};
			{6'd27, 6'd57}: color = {8'd192, 8'd192, 8'd128};
			{6'd28, 6'd57}: color = {8'd128, 8'd128, 8'd64};
			{6'd29, 6'd57}: color = {8'd128, 8'd128, 8'd64};
			{6'd30, 6'd57}: color = {8'd192, 8'd128, 8'd64};
			{6'd31, 6'd57}: color = {8'd192, 8'd128, 8'd128};
			{6'd32, 6'd57}: color = {8'd192, 8'd192, 8'd128};
			{6'd33, 6'd57}: color = {8'd192, 8'd128, 8'd128};
			{6'd34, 6'd57}: color = {8'd192, 8'd128, 8'd64};
			{6'd35, 6'd57}: color = {8'd192, 8'd128, 8'd128};
			{6'd36, 6'd57}: color = {8'd192, 8'd192, 8'd128};
			{6'd37, 6'd57}: color = {8'd192, 8'd128, 8'd128};
			{6'd38, 6'd57}: color = {8'd192, 8'd192, 8'd128};
			{6'd39, 6'd57}: color = {8'd192, 8'd192, 8'd128};
			{6'd40, 6'd57}: color = {8'd192, 8'd128, 8'd64};
			{6'd41, 6'd57}: color = {8'd192, 8'd192, 8'd128};
			{6'd42, 6'd57}: color = {8'd128, 8'd128, 8'd128};
			{6'd43, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd57}: color = {8'd64, 8'd64, 8'd64};
			{6'd47, 6'd57}: color = {8'd128, 8'd128, 8'd128};
			{6'd48, 6'd57}: color = {8'd192, 8'd192, 8'd192};
			{6'd49, 6'd57}: color = {8'd192, 8'd192, 8'd192};
			{6'd50, 6'd57}: color = {8'd192, 8'd192, 8'd192};
			{6'd51, 6'd57}: color = {8'd128, 8'd128, 8'd128};
			{6'd52, 6'd57}: color = {8'd64, 8'd64, 8'd64};
			{6'd53, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd57}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd58}: color = {8'd64, 8'd64, 8'd64};
			{6'd16, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd17, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd18, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd58}: color = {8'd128, 8'd128, 8'd128};
			{6'd21, 6'd58}: color = {8'd64, 8'd64, 8'd64};
			{6'd22, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd27, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd28, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd29, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd30, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd31, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd32, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd33, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd34, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd35, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd36, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd37, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd38, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd39, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd40, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd58}: color = {8'd64, 8'd64, 8'd64};
			{6'd45, 6'd58}: color = {8'd128, 8'd128, 8'd128};
			{6'd46, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd47, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd48, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd49, 6'd58}: color = {8'd192, 8'd192, 8'd192};
			{6'd50, 6'd58}: color = {8'd128, 8'd128, 8'd128};
			{6'd51, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd58}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd59}: color = {8'd64, 8'd64, 8'd64};
			{6'd17, 6'd59}: color = {8'd128, 8'd128, 8'd128};
			{6'd18, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd19, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd20, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd59}: color = {8'd128, 8'd128, 8'd128};
			{6'd23, 6'd59}: color = {8'd128, 8'd128, 8'd128};
			{6'd24, 6'd59}: color = {8'd64, 8'd64, 8'd64};
			{6'd25, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd27, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd28, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd29, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd30, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd31, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd32, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd33, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd34, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd35, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd36, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd37, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd38, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd39, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd40, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd59}: color = {8'd64, 8'd64, 8'd64};
			{6'd42, 6'd59}: color = {8'd128, 8'd128, 8'd128};
			{6'd43, 6'd59}: color = {8'd128, 8'd128, 8'd128};
			{6'd44, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd45, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd46, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd47, 6'd59}: color = {8'd192, 8'd192, 8'd192};
			{6'd48, 6'd59}: color = {8'd128, 8'd128, 8'd128};
			{6'd49, 6'd59}: color = {8'd64, 8'd64, 8'd64};
			{6'd50, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd59}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd19, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd20, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd21, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd22, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd23, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd26, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd27, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd28, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd29, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd30, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd31, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd32, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd33, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd34, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd35, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd36, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd37, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd38, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd39, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd40, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd41, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd42, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd43, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd44, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd45, 6'd60}: color = {8'd192, 8'd192, 8'd192};
			{6'd46, 6'd60}: color = {8'd128, 8'd128, 8'd128};
			{6'd47, 6'd60}: color = {8'd64, 8'd64, 8'd64};
			{6'd48, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd60}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd61}: color = {8'd64, 8'd64, 8'd64};
			{6'd21, 6'd61}: color = {8'd128, 8'd128, 8'd128};
			{6'd22, 6'd61}: color = {8'd128, 8'd128, 8'd128};
			{6'd23, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd24, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd25, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd26, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd32, 6'd61}: color = {8'd128, 8'd128, 8'd128};
			{6'd33, 6'd61}: color = {8'd128, 8'd128, 8'd128};
			{6'd34, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd39, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd40, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd41, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd42, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd43, 6'd61}: color = {8'd192, 8'd192, 8'd192};
			{6'd44, 6'd61}: color = {8'd128, 8'd128, 8'd128};
			{6'd45, 6'd61}: color = {8'd64, 8'd64, 8'd64};
			{6'd46, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd61}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd62}: color = {8'd64, 8'd64, 8'd64};
			{6'd24, 6'd62}: color = {8'd128, 8'd128, 8'd128};
			{6'd25, 6'd62}: color = {8'd128, 8'd128, 8'd128};
			{6'd26, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd27, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd28, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd29, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd30, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd31, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd32, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd33, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd34, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd35, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd36, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd37, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd38, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd39, 6'd62}: color = {8'd192, 8'd192, 8'd192};
			{6'd40, 6'd62}: color = {8'd128, 8'd128, 8'd128};
			{6'd41, 6'd62}: color = {8'd128, 8'd128, 8'd128};
			{6'd42, 6'd62}: color = {8'd64, 8'd64, 8'd64};
			{6'd43, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd62}: color = {8'd0, 8'd0, 8'd0};
			{6'd0, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd1, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd2, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd3, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd4, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd5, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd6, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd7, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd8, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd9, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd10, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd11, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd12, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd13, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd14, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd15, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd16, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd17, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd18, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd19, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd20, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd21, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd22, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd23, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd24, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd25, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd26, 6'd63}: color = {8'd64, 8'd64, 8'd64};
			{6'd27, 6'd63}: color = {8'd64, 8'd64, 8'd64};
			{6'd28, 6'd63}: color = {8'd64, 8'd64, 8'd64};
			{6'd29, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd30, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd31, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd32, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd33, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd34, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd35, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd36, 6'd63}: color = {8'd128, 8'd128, 8'd128};
			{6'd37, 6'd63}: color = {8'd64, 8'd64, 8'd64};
			{6'd38, 6'd63}: color = {8'd64, 8'd64, 8'd64};
			{6'd39, 6'd63}: color = {8'd64, 8'd64, 8'd64};
			{6'd40, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd41, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd42, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd43, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd44, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd45, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd46, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd47, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd48, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd49, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd50, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd51, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd52, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd53, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd54, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd55, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd56, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd57, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd58, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd59, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd60, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd61, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd62, 6'd63}: color = {8'd0, 8'd0, 8'd0};
			{6'd63, 6'd63}: color = {8'd0, 8'd0, 8'd0};
		endcase
endmodule
