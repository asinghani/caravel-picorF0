magic
tech sky130A
magscale 1 2
timestamp 1636925932
<< obsli1 >>
rect 1104 2159 118283 118609
<< obsm1 >>
rect 106 1572 119034 118640
<< metal2 >>
rect 478 120483 534 121283
rect 1490 120483 1546 121283
rect 2502 120483 2558 121283
rect 3606 120483 3662 121283
rect 4618 120483 4674 121283
rect 5630 120483 5686 121283
rect 6734 120483 6790 121283
rect 7746 120483 7802 121283
rect 8758 120483 8814 121283
rect 9862 120483 9918 121283
rect 10874 120483 10930 121283
rect 11886 120483 11942 121283
rect 12990 120483 13046 121283
rect 14002 120483 14058 121283
rect 15106 120483 15162 121283
rect 16118 120483 16174 121283
rect 17130 120483 17186 121283
rect 18234 120483 18290 121283
rect 19246 120483 19302 121283
rect 20258 120483 20314 121283
rect 21362 120483 21418 121283
rect 22374 120483 22430 121283
rect 23386 120483 23442 121283
rect 24490 120483 24546 121283
rect 25502 120483 25558 121283
rect 26514 120483 26570 121283
rect 27618 120483 27674 121283
rect 28630 120483 28686 121283
rect 29734 120483 29790 121283
rect 30746 120483 30802 121283
rect 31758 120483 31814 121283
rect 32862 120483 32918 121283
rect 33874 120483 33930 121283
rect 34886 120483 34942 121283
rect 35990 120483 36046 121283
rect 37002 120483 37058 121283
rect 38014 120483 38070 121283
rect 39118 120483 39174 121283
rect 40130 120483 40186 121283
rect 41234 120483 41290 121283
rect 42246 120483 42302 121283
rect 43258 120483 43314 121283
rect 44362 120483 44418 121283
rect 45374 120483 45430 121283
rect 46386 120483 46442 121283
rect 47490 120483 47546 121283
rect 48502 120483 48558 121283
rect 49514 120483 49570 121283
rect 50618 120483 50674 121283
rect 51630 120483 51686 121283
rect 52642 120483 52698 121283
rect 53746 120483 53802 121283
rect 54758 120483 54814 121283
rect 55862 120483 55918 121283
rect 56874 120483 56930 121283
rect 57886 120483 57942 121283
rect 58990 120483 59046 121283
rect 60002 120483 60058 121283
rect 61014 120483 61070 121283
rect 62118 120483 62174 121283
rect 63130 120483 63186 121283
rect 64142 120483 64198 121283
rect 65246 120483 65302 121283
rect 66258 120483 66314 121283
rect 67362 120483 67418 121283
rect 68374 120483 68430 121283
rect 69386 120483 69442 121283
rect 70490 120483 70546 121283
rect 71502 120483 71558 121283
rect 72514 120483 72570 121283
rect 73618 120483 73674 121283
rect 74630 120483 74686 121283
rect 75642 120483 75698 121283
rect 76746 120483 76802 121283
rect 77758 120483 77814 121283
rect 78770 120483 78826 121283
rect 79874 120483 79930 121283
rect 80886 120483 80942 121283
rect 81990 120483 82046 121283
rect 83002 120483 83058 121283
rect 84014 120483 84070 121283
rect 85118 120483 85174 121283
rect 86130 120483 86186 121283
rect 87142 120483 87198 121283
rect 88246 120483 88302 121283
rect 89258 120483 89314 121283
rect 90270 120483 90326 121283
rect 91374 120483 91430 121283
rect 92386 120483 92442 121283
rect 93490 120483 93546 121283
rect 94502 120483 94558 121283
rect 95514 120483 95570 121283
rect 96618 120483 96674 121283
rect 97630 120483 97686 121283
rect 98642 120483 98698 121283
rect 99746 120483 99802 121283
rect 100758 120483 100814 121283
rect 101770 120483 101826 121283
rect 102874 120483 102930 121283
rect 103886 120483 103942 121283
rect 104898 120483 104954 121283
rect 106002 120483 106058 121283
rect 107014 120483 107070 121283
rect 108118 120483 108174 121283
rect 109130 120483 109186 121283
rect 110142 120483 110198 121283
rect 111246 120483 111302 121283
rect 112258 120483 112314 121283
rect 113270 120483 113326 121283
rect 114374 120483 114430 121283
rect 115386 120483 115442 121283
rect 116398 120483 116454 121283
rect 117502 120483 117558 121283
rect 118514 120483 118570 121283
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3422 0 3478 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7102 0 7158 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39210 0 39266 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47674 0 47730 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51538 0 51594 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 53010 0 53066 800
rect 53194 0 53250 800
rect 53470 0 53526 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56138 0 56194 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61934 0 61990 800
rect 62210 0 62266 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65798 0 65854 800
rect 66074 0 66130 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77666 0 77722 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78586 0 78642 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81530 0 81586 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82266 0 82322 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86590 0 86646 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87786 0 87842 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89258 0 89314 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 89994 0 90050 800
rect 90178 0 90234 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96986 0 97042 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 97906 0 97962 800
rect 98182 0 98238 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100574 0 100630 800
rect 100850 0 100906 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101586 0 101642 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102322 0 102378 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103242 0 103298 800
rect 103518 0 103574 800
rect 103702 0 103758 800
rect 103978 0 104034 800
rect 104254 0 104310 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105174 0 105230 800
rect 105450 0 105506 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106370 0 106426 800
rect 106646 0 106702 800
rect 106922 0 106978 800
rect 107106 0 107162 800
rect 107382 0 107438 800
rect 107566 0 107622 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108302 0 108358 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109038 0 109094 800
rect 109314 0 109370 800
rect 109498 0 109554 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110786 0 110842 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111430 0 111486 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112166 0 112222 800
rect 112442 0 112498 800
rect 112718 0 112774 800
rect 112902 0 112958 800
rect 113178 0 113234 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114098 0 114154 800
rect 114374 0 114430 800
rect 114650 0 114706 800
rect 114834 0 114890 800
rect 115110 0 115166 800
rect 115294 0 115350 800
rect 115570 0 115626 800
rect 115846 0 115902 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116766 0 116822 800
rect 117042 0 117098 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 117962 0 118018 800
rect 118238 0 118294 800
rect 118514 0 118570 800
rect 118698 0 118754 800
rect 118974 0 119030 800
<< obsm2 >>
rect 112 120427 422 120483
rect 590 120427 1434 120483
rect 1602 120427 2446 120483
rect 2614 120427 3550 120483
rect 3718 120427 4562 120483
rect 4730 120427 5574 120483
rect 5742 120427 6678 120483
rect 6846 120427 7690 120483
rect 7858 120427 8702 120483
rect 8870 120427 9806 120483
rect 9974 120427 10818 120483
rect 10986 120427 11830 120483
rect 11998 120427 12934 120483
rect 13102 120427 13946 120483
rect 14114 120427 15050 120483
rect 15218 120427 16062 120483
rect 16230 120427 17074 120483
rect 17242 120427 18178 120483
rect 18346 120427 19190 120483
rect 19358 120427 20202 120483
rect 20370 120427 21306 120483
rect 21474 120427 22318 120483
rect 22486 120427 23330 120483
rect 23498 120427 24434 120483
rect 24602 120427 25446 120483
rect 25614 120427 26458 120483
rect 26626 120427 27562 120483
rect 27730 120427 28574 120483
rect 28742 120427 29678 120483
rect 29846 120427 30690 120483
rect 30858 120427 31702 120483
rect 31870 120427 32806 120483
rect 32974 120427 33818 120483
rect 33986 120427 34830 120483
rect 34998 120427 35934 120483
rect 36102 120427 36946 120483
rect 37114 120427 37958 120483
rect 38126 120427 39062 120483
rect 39230 120427 40074 120483
rect 40242 120427 41178 120483
rect 41346 120427 42190 120483
rect 42358 120427 43202 120483
rect 43370 120427 44306 120483
rect 44474 120427 45318 120483
rect 45486 120427 46330 120483
rect 46498 120427 47434 120483
rect 47602 120427 48446 120483
rect 48614 120427 49458 120483
rect 49626 120427 50562 120483
rect 50730 120427 51574 120483
rect 51742 120427 52586 120483
rect 52754 120427 53690 120483
rect 53858 120427 54702 120483
rect 54870 120427 55806 120483
rect 55974 120427 56818 120483
rect 56986 120427 57830 120483
rect 57998 120427 58934 120483
rect 59102 120427 59946 120483
rect 60114 120427 60958 120483
rect 61126 120427 62062 120483
rect 62230 120427 63074 120483
rect 63242 120427 64086 120483
rect 64254 120427 65190 120483
rect 65358 120427 66202 120483
rect 66370 120427 67306 120483
rect 67474 120427 68318 120483
rect 68486 120427 69330 120483
rect 69498 120427 70434 120483
rect 70602 120427 71446 120483
rect 71614 120427 72458 120483
rect 72626 120427 73562 120483
rect 73730 120427 74574 120483
rect 74742 120427 75586 120483
rect 75754 120427 76690 120483
rect 76858 120427 77702 120483
rect 77870 120427 78714 120483
rect 78882 120427 79818 120483
rect 79986 120427 80830 120483
rect 80998 120427 81934 120483
rect 82102 120427 82946 120483
rect 83114 120427 83958 120483
rect 84126 120427 85062 120483
rect 85230 120427 86074 120483
rect 86242 120427 87086 120483
rect 87254 120427 88190 120483
rect 88358 120427 89202 120483
rect 89370 120427 90214 120483
rect 90382 120427 91318 120483
rect 91486 120427 92330 120483
rect 92498 120427 93434 120483
rect 93602 120427 94446 120483
rect 94614 120427 95458 120483
rect 95626 120427 96562 120483
rect 96730 120427 97574 120483
rect 97742 120427 98586 120483
rect 98754 120427 99690 120483
rect 99858 120427 100702 120483
rect 100870 120427 101714 120483
rect 101882 120427 102818 120483
rect 102986 120427 103830 120483
rect 103998 120427 104842 120483
rect 105010 120427 105946 120483
rect 106114 120427 106958 120483
rect 107126 120427 108062 120483
rect 108230 120427 109074 120483
rect 109242 120427 110086 120483
rect 110254 120427 111190 120483
rect 111358 120427 112202 120483
rect 112370 120427 113214 120483
rect 113382 120427 114318 120483
rect 114486 120427 115330 120483
rect 115498 120427 116342 120483
rect 116510 120427 117446 120483
rect 117614 120427 118458 120483
rect 118626 120427 119028 120483
rect 112 856 119028 120427
rect 222 800 238 856
rect 406 800 514 856
rect 682 800 698 856
rect 866 800 974 856
rect 1142 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1710 856
rect 1878 800 1986 856
rect 2154 800 2170 856
rect 2338 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2906 856
rect 3074 800 3182 856
rect 3350 800 3366 856
rect 3534 800 3642 856
rect 3810 800 3918 856
rect 4086 800 4102 856
rect 4270 800 4378 856
rect 4546 800 4562 856
rect 4730 800 4838 856
rect 5006 800 5114 856
rect 5282 800 5298 856
rect 5466 800 5574 856
rect 5742 800 5850 856
rect 6018 800 6034 856
rect 6202 800 6310 856
rect 6478 800 6494 856
rect 6662 800 6770 856
rect 6938 800 7046 856
rect 7214 800 7230 856
rect 7398 800 7506 856
rect 7674 800 7782 856
rect 7950 800 7966 856
rect 8134 800 8242 856
rect 8410 800 8426 856
rect 8594 800 8702 856
rect 8870 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9438 856
rect 9606 800 9714 856
rect 9882 800 9898 856
rect 10066 800 10174 856
rect 10342 800 10358 856
rect 10526 800 10634 856
rect 10802 800 10910 856
rect 11078 800 11094 856
rect 11262 800 11370 856
rect 11538 800 11646 856
rect 11814 800 11830 856
rect 11998 800 12106 856
rect 12274 800 12290 856
rect 12458 800 12566 856
rect 12734 800 12842 856
rect 13010 800 13026 856
rect 13194 800 13302 856
rect 13470 800 13578 856
rect 13746 800 13762 856
rect 13930 800 14038 856
rect 14206 800 14222 856
rect 14390 800 14498 856
rect 14666 800 14774 856
rect 14942 800 14958 856
rect 15126 800 15234 856
rect 15402 800 15510 856
rect 15678 800 15694 856
rect 15862 800 15970 856
rect 16138 800 16154 856
rect 16322 800 16430 856
rect 16598 800 16706 856
rect 16874 800 16890 856
rect 17058 800 17166 856
rect 17334 800 17442 856
rect 17610 800 17626 856
rect 17794 800 17902 856
rect 18070 800 18178 856
rect 18346 800 18362 856
rect 18530 800 18638 856
rect 18806 800 18822 856
rect 18990 800 19098 856
rect 19266 800 19374 856
rect 19542 800 19558 856
rect 19726 800 19834 856
rect 20002 800 20110 856
rect 20278 800 20294 856
rect 20462 800 20570 856
rect 20738 800 20754 856
rect 20922 800 21030 856
rect 21198 800 21306 856
rect 21474 800 21490 856
rect 21658 800 21766 856
rect 21934 800 22042 856
rect 22210 800 22226 856
rect 22394 800 22502 856
rect 22670 800 22686 856
rect 22854 800 22962 856
rect 23130 800 23238 856
rect 23406 800 23422 856
rect 23590 800 23698 856
rect 23866 800 23974 856
rect 24142 800 24158 856
rect 24326 800 24434 856
rect 24602 800 24618 856
rect 24786 800 24894 856
rect 25062 800 25170 856
rect 25338 800 25354 856
rect 25522 800 25630 856
rect 25798 800 25906 856
rect 26074 800 26090 856
rect 26258 800 26366 856
rect 26534 800 26550 856
rect 26718 800 26826 856
rect 26994 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27562 856
rect 27730 800 27838 856
rect 28006 800 28022 856
rect 28190 800 28298 856
rect 28466 800 28482 856
rect 28650 800 28758 856
rect 28926 800 29034 856
rect 29202 800 29218 856
rect 29386 800 29494 856
rect 29662 800 29770 856
rect 29938 800 29954 856
rect 30122 800 30230 856
rect 30398 800 30414 856
rect 30582 800 30690 856
rect 30858 800 30966 856
rect 31134 800 31150 856
rect 31318 800 31426 856
rect 31594 800 31702 856
rect 31870 800 31886 856
rect 32054 800 32162 856
rect 32330 800 32346 856
rect 32514 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33082 856
rect 33250 800 33358 856
rect 33526 800 33634 856
rect 33802 800 33818 856
rect 33986 800 34094 856
rect 34262 800 34370 856
rect 34538 800 34554 856
rect 34722 800 34830 856
rect 34998 800 35014 856
rect 35182 800 35290 856
rect 35458 800 35566 856
rect 35734 800 35750 856
rect 35918 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36762 856
rect 36930 800 36946 856
rect 37114 800 37222 856
rect 37390 800 37498 856
rect 37666 800 37682 856
rect 37850 800 37958 856
rect 38126 800 38234 856
rect 38402 800 38418 856
rect 38586 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39154 856
rect 39322 800 39430 856
rect 39598 800 39614 856
rect 39782 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40626 856
rect 40794 800 40810 856
rect 40978 800 41086 856
rect 41254 800 41362 856
rect 41530 800 41546 856
rect 41714 800 41822 856
rect 41990 800 42098 856
rect 42266 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42742 856
rect 42910 800 43018 856
rect 43186 800 43294 856
rect 43462 800 43478 856
rect 43646 800 43754 856
rect 43922 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44674 856
rect 44842 800 44950 856
rect 45118 800 45226 856
rect 45394 800 45410 856
rect 45578 800 45686 856
rect 45854 800 45962 856
rect 46130 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46882 856
rect 47050 800 47158 856
rect 47326 800 47342 856
rect 47510 800 47618 856
rect 47786 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48354 856
rect 48522 800 48538 856
rect 48706 800 48814 856
rect 48982 800 49090 856
rect 49258 800 49274 856
rect 49442 800 49550 856
rect 49718 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50286 856
rect 50454 800 50470 856
rect 50638 800 50746 856
rect 50914 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51482 856
rect 51650 800 51758 856
rect 51926 800 51942 856
rect 52110 800 52218 856
rect 52386 800 52494 856
rect 52662 800 52678 856
rect 52846 800 52954 856
rect 53122 800 53138 856
rect 53306 800 53414 856
rect 53582 800 53690 856
rect 53858 800 53874 856
rect 54042 800 54150 856
rect 54318 800 54426 856
rect 54594 800 54610 856
rect 54778 800 54886 856
rect 55054 800 55070 856
rect 55238 800 55346 856
rect 55514 800 55622 856
rect 55790 800 55806 856
rect 55974 800 56082 856
rect 56250 800 56358 856
rect 56526 800 56542 856
rect 56710 800 56818 856
rect 56986 800 57002 856
rect 57170 800 57278 856
rect 57446 800 57554 856
rect 57722 800 57738 856
rect 57906 800 58014 856
rect 58182 800 58290 856
rect 58458 800 58474 856
rect 58642 800 58750 856
rect 58918 800 58934 856
rect 59102 800 59210 856
rect 59378 800 59486 856
rect 59654 800 59670 856
rect 59838 800 59946 856
rect 60114 800 60222 856
rect 60390 800 60406 856
rect 60574 800 60682 856
rect 60850 800 60866 856
rect 61034 800 61142 856
rect 61310 800 61418 856
rect 61586 800 61602 856
rect 61770 800 61878 856
rect 62046 800 62154 856
rect 62322 800 62338 856
rect 62506 800 62614 856
rect 62782 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63350 856
rect 63518 800 63534 856
rect 63702 800 63810 856
rect 63978 800 64086 856
rect 64254 800 64270 856
rect 64438 800 64546 856
rect 64714 800 64730 856
rect 64898 800 65006 856
rect 65174 800 65282 856
rect 65450 800 65466 856
rect 65634 800 65742 856
rect 65910 800 66018 856
rect 66186 800 66202 856
rect 66370 800 66478 856
rect 66646 800 66662 856
rect 66830 800 66938 856
rect 67106 800 67214 856
rect 67382 800 67398 856
rect 67566 800 67674 856
rect 67842 800 67950 856
rect 68118 800 68134 856
rect 68302 800 68410 856
rect 68578 800 68686 856
rect 68854 800 68870 856
rect 69038 800 69146 856
rect 69314 800 69330 856
rect 69498 800 69606 856
rect 69774 800 69882 856
rect 70050 800 70066 856
rect 70234 800 70342 856
rect 70510 800 70618 856
rect 70786 800 70802 856
rect 70970 800 71078 856
rect 71246 800 71262 856
rect 71430 800 71538 856
rect 71706 800 71814 856
rect 71982 800 71998 856
rect 72166 800 72274 856
rect 72442 800 72550 856
rect 72718 800 72734 856
rect 72902 800 73010 856
rect 73178 800 73194 856
rect 73362 800 73470 856
rect 73638 800 73746 856
rect 73914 800 73930 856
rect 74098 800 74206 856
rect 74374 800 74482 856
rect 74650 800 74666 856
rect 74834 800 74942 856
rect 75110 800 75126 856
rect 75294 800 75402 856
rect 75570 800 75678 856
rect 75846 800 75862 856
rect 76030 800 76138 856
rect 76306 800 76414 856
rect 76582 800 76598 856
rect 76766 800 76874 856
rect 77042 800 77058 856
rect 77226 800 77334 856
rect 77502 800 77610 856
rect 77778 800 77794 856
rect 77962 800 78070 856
rect 78238 800 78346 856
rect 78514 800 78530 856
rect 78698 800 78806 856
rect 78974 800 78990 856
rect 79158 800 79266 856
rect 79434 800 79542 856
rect 79710 800 79726 856
rect 79894 800 80002 856
rect 80170 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80738 856
rect 80906 800 80922 856
rect 81090 800 81198 856
rect 81366 800 81474 856
rect 81642 800 81658 856
rect 81826 800 81934 856
rect 82102 800 82210 856
rect 82378 800 82394 856
rect 82562 800 82670 856
rect 82838 800 82854 856
rect 83022 800 83130 856
rect 83298 800 83406 856
rect 83574 800 83590 856
rect 83758 800 83866 856
rect 84034 800 84142 856
rect 84310 800 84326 856
rect 84494 800 84602 856
rect 84770 800 84786 856
rect 84954 800 85062 856
rect 85230 800 85338 856
rect 85506 800 85522 856
rect 85690 800 85798 856
rect 85966 800 86074 856
rect 86242 800 86258 856
rect 86426 800 86534 856
rect 86702 800 86810 856
rect 86978 800 86994 856
rect 87162 800 87270 856
rect 87438 800 87454 856
rect 87622 800 87730 856
rect 87898 800 88006 856
rect 88174 800 88190 856
rect 88358 800 88466 856
rect 88634 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89202 856
rect 89370 800 89386 856
rect 89554 800 89662 856
rect 89830 800 89938 856
rect 90106 800 90122 856
rect 90290 800 90398 856
rect 90566 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91134 856
rect 91302 800 91318 856
rect 91486 800 91594 856
rect 91762 800 91870 856
rect 92038 800 92054 856
rect 92222 800 92330 856
rect 92498 800 92606 856
rect 92774 800 92790 856
rect 92958 800 93066 856
rect 93234 800 93250 856
rect 93418 800 93526 856
rect 93694 800 93802 856
rect 93970 800 93986 856
rect 94154 800 94262 856
rect 94430 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94998 856
rect 95166 800 95182 856
rect 95350 800 95458 856
rect 95626 800 95734 856
rect 95902 800 95918 856
rect 96086 800 96194 856
rect 96362 800 96470 856
rect 96638 800 96654 856
rect 96822 800 96930 856
rect 97098 800 97114 856
rect 97282 800 97390 856
rect 97558 800 97666 856
rect 97834 800 97850 856
rect 98018 800 98126 856
rect 98294 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98862 856
rect 99030 800 99046 856
rect 99214 800 99322 856
rect 99490 800 99598 856
rect 99766 800 99782 856
rect 99950 800 100058 856
rect 100226 800 100334 856
rect 100502 800 100518 856
rect 100686 800 100794 856
rect 100962 800 100978 856
rect 101146 800 101254 856
rect 101422 800 101530 856
rect 101698 800 101714 856
rect 101882 800 101990 856
rect 102158 800 102266 856
rect 102434 800 102450 856
rect 102618 800 102726 856
rect 102894 800 103002 856
rect 103170 800 103186 856
rect 103354 800 103462 856
rect 103630 800 103646 856
rect 103814 800 103922 856
rect 104090 800 104198 856
rect 104366 800 104382 856
rect 104550 800 104658 856
rect 104826 800 104934 856
rect 105102 800 105118 856
rect 105286 800 105394 856
rect 105562 800 105578 856
rect 105746 800 105854 856
rect 106022 800 106130 856
rect 106298 800 106314 856
rect 106482 800 106590 856
rect 106758 800 106866 856
rect 107034 800 107050 856
rect 107218 800 107326 856
rect 107494 800 107510 856
rect 107678 800 107786 856
rect 107954 800 108062 856
rect 108230 800 108246 856
rect 108414 800 108522 856
rect 108690 800 108798 856
rect 108966 800 108982 856
rect 109150 800 109258 856
rect 109426 800 109442 856
rect 109610 800 109718 856
rect 109886 800 109994 856
rect 110162 800 110178 856
rect 110346 800 110454 856
rect 110622 800 110730 856
rect 110898 800 110914 856
rect 111082 800 111190 856
rect 111358 800 111374 856
rect 111542 800 111650 856
rect 111818 800 111926 856
rect 112094 800 112110 856
rect 112278 800 112386 856
rect 112554 800 112662 856
rect 112830 800 112846 856
rect 113014 800 113122 856
rect 113290 800 113306 856
rect 113474 800 113582 856
rect 113750 800 113858 856
rect 114026 800 114042 856
rect 114210 800 114318 856
rect 114486 800 114594 856
rect 114762 800 114778 856
rect 114946 800 115054 856
rect 115222 800 115238 856
rect 115406 800 115514 856
rect 115682 800 115790 856
rect 115958 800 115974 856
rect 116142 800 116250 856
rect 116418 800 116526 856
rect 116694 800 116710 856
rect 116878 800 116986 856
rect 117154 800 117170 856
rect 117338 800 117446 856
rect 117614 800 117722 856
rect 117890 800 117906 856
rect 118074 800 118182 856
rect 118350 800 118458 856
rect 118626 800 118642 856
rect 118810 800 118918 856
<< obsm3 >>
rect 3049 2143 113423 118625
<< metal4 >>
rect 4208 2128 4528 118640
rect 19568 2128 19888 118640
rect 34928 2128 35248 118640
rect 50288 2128 50608 118640
rect 65648 2128 65968 118640
rect 81008 2128 81328 118640
rect 96368 2128 96688 118640
rect 111728 2128 112048 118640
<< obsm4 >>
rect 4843 55931 19488 115429
rect 19968 55931 34848 115429
rect 35328 55931 50208 115429
rect 50688 55931 65568 115429
rect 66048 55931 69309 115429
<< labels >>
rlabel metal2 s 478 120483 534 121283 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 31758 120483 31814 121283 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 34886 120483 34942 121283 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 38014 120483 38070 121283 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 41234 120483 41290 121283 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 44362 120483 44418 121283 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 47490 120483 47546 121283 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 50618 120483 50674 121283 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 53746 120483 53802 121283 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 56874 120483 56930 121283 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 60002 120483 60058 121283 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3606 120483 3662 121283 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 63130 120483 63186 121283 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 66258 120483 66314 121283 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 69386 120483 69442 121283 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 72514 120483 72570 121283 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 75642 120483 75698 121283 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 78770 120483 78826 121283 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 81990 120483 82046 121283 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 85118 120483 85174 121283 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 88246 120483 88302 121283 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 91374 120483 91430 121283 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6734 120483 6790 121283 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 94502 120483 94558 121283 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 97630 120483 97686 121283 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 100758 120483 100814 121283 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 103886 120483 103942 121283 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 107014 120483 107070 121283 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 110142 120483 110198 121283 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 113270 120483 113326 121283 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 116398 120483 116454 121283 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9862 120483 9918 121283 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12990 120483 13046 121283 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 16118 120483 16174 121283 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 19246 120483 19302 121283 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 22374 120483 22430 121283 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 25502 120483 25558 121283 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 28630 120483 28686 121283 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1490 120483 1546 121283 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 32862 120483 32918 121283 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 35990 120483 36046 121283 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 39118 120483 39174 121283 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 42246 120483 42302 121283 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 45374 120483 45430 121283 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 48502 120483 48558 121283 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 51630 120483 51686 121283 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 54758 120483 54814 121283 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 57886 120483 57942 121283 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 61014 120483 61070 121283 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4618 120483 4674 121283 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 64142 120483 64198 121283 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 67362 120483 67418 121283 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 70490 120483 70546 121283 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 73618 120483 73674 121283 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 76746 120483 76802 121283 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 79874 120483 79930 121283 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 83002 120483 83058 121283 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 86130 120483 86186 121283 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 89258 120483 89314 121283 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 92386 120483 92442 121283 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7746 120483 7802 121283 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 95514 120483 95570 121283 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 98642 120483 98698 121283 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 101770 120483 101826 121283 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 104898 120483 104954 121283 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 108118 120483 108174 121283 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 111246 120483 111302 121283 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 114374 120483 114430 121283 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 117502 120483 117558 121283 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10874 120483 10930 121283 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 14002 120483 14058 121283 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 17130 120483 17186 121283 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 20258 120483 20314 121283 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 23386 120483 23442 121283 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 26514 120483 26570 121283 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 29734 120483 29790 121283 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2502 120483 2558 121283 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 33874 120483 33930 121283 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 37002 120483 37058 121283 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 40130 120483 40186 121283 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 43258 120483 43314 121283 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 46386 120483 46442 121283 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 49514 120483 49570 121283 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 52642 120483 52698 121283 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 55862 120483 55918 121283 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 58990 120483 59046 121283 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 62118 120483 62174 121283 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5630 120483 5686 121283 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 65246 120483 65302 121283 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 68374 120483 68430 121283 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 71502 120483 71558 121283 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 74630 120483 74686 121283 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 77758 120483 77814 121283 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 80886 120483 80942 121283 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 84014 120483 84070 121283 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 87142 120483 87198 121283 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 90270 120483 90326 121283 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 93490 120483 93546 121283 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8758 120483 8814 121283 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 96618 120483 96674 121283 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 99746 120483 99802 121283 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 102874 120483 102930 121283 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 106002 120483 106058 121283 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 109130 120483 109186 121283 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 112258 120483 112314 121283 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 115386 120483 115442 121283 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 118514 120483 118570 121283 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11886 120483 11942 121283 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 15106 120483 15162 121283 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 18234 120483 18290 121283 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 21362 120483 21418 121283 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 24490 120483 24546 121283 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 27618 120483 27674 121283 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 30746 120483 30802 121283 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 118974 0 119030 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 118640 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 118640 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 118640 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 118640 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 118640 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 118640 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 118640 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 118640 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 119139 121283
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 27905838
string GDS_START 1194960
<< end >>

