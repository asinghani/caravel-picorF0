// SPDX-FileCopyrightText: 2021 Natalia Machado
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype wire
/* Generated by Yosys 0.11 (git sha1 UNKNOWN, clang 10.0.1 -fPIC -Os) */
(* cells_not_processed =  1  *)
module CanAcf(clock, reset, io_id, io_resetMode, io_acceptanceFilterMode, io_extendedMode, io_acceptanceCode_0, io_acceptanceCode_1, io_acceptanceCode_2, io_acceptanceCode_3, io_acceptanceMask_0, io_acceptanceMask_1, io_acceptanceMask_2, io_acceptanceMask_3, io_goRxCrcLim, io_goRxInter, io_goErrorFrame, io_data0, io_data1, io_rtr1, io_rtr2
, io_ide, io_noByte0, io_noByte1, io_idOk);
  (* src = "CanAcf.scala:60.61|CanAcf.scala:61.10|CanAcf.scala:27.28" *)
  wire _000_;
  (* src = "CanAcf.scala:58.23|CanAcf.scala:59.10" *)
  wire _001_;
  (* src = "CanAcf.scala:60.27" *)
  wire _002_;
  (* src = "CanAcf.scala:60.42" *)
  wire _003_;
  (* src = "CanAcf.scala:33.43" *)
  wire [7:0] _004_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _005_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _006_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _007_;
  (* src = "CanAcf.scala:59.64" *)
  wire _008_;
  (* src = "CanAcf.scala:59.98" *)
  wire _009_;
  (* src = "CanAcf.scala:59.36" *)
  wire _010_;
  (* src = "CanAcf.scala:59.16" *)
  wire _011_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _012_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _013_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _014_;
  (* src = "CanAcf.scala:31.35" *)
  wire _015_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _016_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _017_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _018_;
  (* src = "CanAcf.scala:31.35" *)
  wire _019_;
  (* src = "CanAcf.scala:55.92" *)
  wire _020_;
  (* src = "CanAcf.scala:48.53" *)
  wire [3:0] _021_;
  (* src = "CanAcf.scala:48.80" *)
  wire [3:0] _022_;
  (* src = "CanAcf.scala:31.11" *)
  wire [3:0] _023_;
  (* src = "CanAcf.scala:31.7" *)
  wire [3:0] _024_;
  (* src = "CanAcf.scala:31.26" *)
  wire [3:0] _025_;
  (* src = "CanAcf.scala:31.35" *)
  wire _026_;
  (* src = "CanAcf.scala:48.87" *)
  wire _027_;
  (* src = "CanAcf.scala:47.94" *)
  wire _028_;
  (* src = "CanAcf.scala:49.26" *)
  wire [3:0] _029_;
  (* src = "CanAcf.scala:49.53" *)
  wire [3:0] _030_;
  (* src = "CanAcf.scala:49.80" *)
  wire [3:0] _031_;
  (* src = "CanAcf.scala:31.11" *)
  wire [3:0] _032_;
  (* src = "CanAcf.scala:31.7" *)
  wire [3:0] _033_;
  (* src = "CanAcf.scala:31.26" *)
  wire [3:0] _034_;
  (* src = "CanAcf.scala:31.35" *)
  wire _035_;
  (* src = "CanAcf.scala:49.87" *)
  wire _036_;
  (* src = "CanAcf.scala:48.101" *)
  wire _037_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _038_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _039_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _040_;
  (* src = "CanAcf.scala:31.35" *)
  wire _041_;
  (* src = "CanAcf.scala:51.61" *)
  wire [3:0] _042_;
  (* src = "CanAcf.scala:51.87" *)
  wire [3:0] _043_;
  (* src = "CanAcf.scala:31.11" *)
  wire [3:0] _044_;
  (* src = "CanAcf.scala:31.7" *)
  wire [3:0] _045_;
  (* src = "CanAcf.scala:31.26" *)
  wire [3:0] _046_;
  (* src = "CanAcf.scala:31.35" *)
  wire _047_;
  (* src = "CanAcf.scala:50.75" *)
  wire _048_;
  (* src = "CanAcf.scala:48.26" *)
  wire [3:0] _049_;
  (* src = "CanAcf.scala:40.44" *)
  wire [7:0] _050_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _051_;
  (* src = "CanAcf.scala:40.97" *)
  wire _052_;
  (* src = "CanAcf.scala:42.22" *)
  wire [7:0] _053_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _054_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _055_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _056_;
  (* src = "CanAcf.scala:31.35" *)
  wire _057_;
  (* src = "CanAcf.scala:41.75" *)
  wire _058_;
  (* src = "CanAcf.scala:43.26" *)
  wire [4:0] _059_;
  (* src = "Cat.scala:30.58" *)
  wire [5:0] _060_;
  (* src = "CanAcf.scala:43.61" *)
  wire [5:0] _061_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _062_;
  (* src = "CanAcf.scala:43.87" *)
  wire [5:0] _063_;
  (* src = "CanAcf.scala:31.11" *)
  wire [5:0] _064_;
  (* src = "CanAcf.scala:31.7" *)
  wire [5:0] _065_;
  (* src = "CanAcf.scala:31.26" *)
  wire [5:0] _066_;
  (* src = "CanAcf.scala:31.35" *)
  wire _067_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _068_;
  (* src = "CanAcf.scala:31.35" *)
  wire _069_;
  (* src = "CanAcf.scala:41.22" *)
  wire [7:0] _070_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _071_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _072_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _073_;
  (* src = "CanAcf.scala:31.35" *)
  wire _074_;
  (* src = "CanAcf.scala:36.26" *)
  wire [2:0] _075_;
  (* src = "Cat.scala:30.58" *)
  wire [3:0] _076_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _077_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _078_;
  (* src = "CanAcf.scala:31.35" *)
  wire _079_;
  (* src = "CanAcf.scala:37.72" *)
  wire _080_;
  (* src = "CanAcf.scala:36.95" *)
  wire _081_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _082_;
  (* src = "CanAcf.scala:31.7" *)
  wire [7:0] _083_;
  (* src = "CanAcf.scala:31.26" *)
  wire [7:0] _084_;
  (* src = "CanAcf.scala:31.35" *)
  wire _085_;
  (* src = "CanAcf.scala:38.72" *)
  wire _086_;
  (* src = "CanAcf.scala:36.61" *)
  wire [3:0] _087_;
  (* src = "CanAcf.scala:36.88" *)
  wire [3:0] _088_;
  (* src = "CanAcf.scala:31.11" *)
  wire [3:0] _089_;
  (* src = "CanAcf.scala:31.7" *)
  wire [3:0] _090_;
  (* src = "CanAcf.scala:31.26" *)
  wire [3:0] _091_;
  (* src = "CanAcf.scala:31.35" *)
  wire _092_;
  (* src = "CanAcf.scala:35.35" *)
  wire _093_;
  (* src = "CanAcf.scala:31.11" *)
  wire [7:0] _094_;
  wire _095_;
  wire _096_;
  input clock;
  (* src = "CanAcf.scala:31.35" *)
  wire idMatch;
  (* src = "CanAcf.scala:27.28" *)
  reg idOk;
  (* src = "CanAcf.scala:27.28|CanAcf.scala:27.28" *)
  wire \idOk$process$CanAcf ;
  input [7:0] io_acceptanceCode_0;
  input [7:0] io_acceptanceCode_1;
  input [7:0] io_acceptanceCode_2;
  input [7:0] io_acceptanceCode_3;
  input io_acceptanceFilterMode;
  input [7:0] io_acceptanceMask_0;
  input [7:0] io_acceptanceMask_1;
  input [7:0] io_acceptanceMask_2;
  input [7:0] io_acceptanceMask_3;
  input [7:0] io_data0;
  input [7:0] io_data1;
  input io_extendedMode;
  input io_goErrorFrame;
  input io_goRxCrcLim;
  input io_goRxInter;
  input [28:0] io_id;
  output io_idOk;
  input io_ide;
  input io_noByte0;
  input io_noByte1;
  input io_resetMode;
  input io_rtr1;
  input io_rtr2;
  (* src = "CanAcf.scala:54.93" *)
  wire matchDfExt;
  (* src = "CanAcf.scala:49.102" *)
  wire matchDfStd;
  (* src = "CanAcf.scala:42.74" *)
  wire matchSfExt;
  (* src = "CanAcf.scala:37.86" *)
  wire matchSfStd;
  input reset;
  assign _093_ = idMatch & _092_;
  assign _081_ = _093_ & _080_;
  assign matchSfStd = _081_ & _086_;
  assign _052_ = _069_ & _074_;
  assign _058_ = _052_ & _057_;
  assign matchSfExt = _058_ & _067_;
  assign _028_ = _093_ & _027_;
  assign _037_ = _028_ & _036_;
  assign _048_ = _041_ & _047_;
  assign _020_ = _015_ & _019_;
  assign _008_ = io_ide ? (* src = "CanAcf.scala:59.64" *) matchSfExt : matchSfStd;
  assign _009_ = io_ide ? (* src = "CanAcf.scala:59.98" *) matchDfExt : matchDfStd;
  assign _010_ = io_acceptanceFilterMode ? (* src = "CanAcf.scala:59.36" *) _008_ : _009_;
  assign _011_ = io_extendedMode ? (* src = "CanAcf.scala:59.16" *) _010_ : idMatch;
  assign _000_ = _003_ ? (* src = "CanAcf.scala:60.61|CanAcf.scala:61.10|CanAcf.scala:27.28" *) 1'h0 : idOk;
  assign _001_ = io_goRxCrcLim ? (* src = "CanAcf.scala:58.23|CanAcf.scala:59.10" *) _011_ : _000_;
  assign _006_ = ~ _005_;
  assign _090_ = ~ _089_;
  assign _077_ = ~ _094_;
  assign _045_ = ~ _044_;
  assign _013_ = ~ _012_;
  assign _017_ = ~ _016_;
  assign _083_ = ~ _082_;
  assign _062_ = ~ _051_;
  assign _072_ = ~ _071_;
  assign _055_ = ~ _054_;
  assign _065_ = ~ _064_;
  assign _024_ = ~ _023_;
  assign _033_ = ~ _032_;
  assign _039_ = ~ _038_;
  assign _007_ = _006_ | io_acceptanceMask_0;
  assign _091_ = _090_ | _088_;
  assign _078_ = _077_ | io_acceptanceMask_2;
  assign _027_ = _026_ | io_noByte0;
  assign _034_ = _033_ | _031_;
  assign _036_ = _035_ | io_noByte0;
  assign _040_ = _039_ | io_acceptanceMask_2;
  assign _046_ = _045_ | _043_;
  assign matchDfStd = _037_ | _048_;
  assign _014_ = _013_ | io_acceptanceMask_2;
  assign _018_ = _017_ | io_acceptanceMask_3;
  assign matchDfExt = _052_ | _020_;
  assign _002_ = io_resetMode | io_goRxInter;
  assign _080_ = _079_ | io_noByte0;
  assign _003_ = _002_ | io_goErrorFrame;
  assign _084_ = _083_ | io_acceptanceMask_3;
  assign _086_ = _085_ | io_noByte1;
  assign _068_ = _062_ | io_acceptanceMask_0;
  assign _073_ = _072_ | io_acceptanceMask_1;
  assign _056_ = _055_ | io_acceptanceMask_2;
  assign _066_ = _065_ | _063_;
  assign _025_ = _024_ | _022_;
  always @(posedge clock)
    idOk <= _095_;
  assign _095_ = _096_ ? (* full_case = 32'd1 *) (* src = "CanAcf.scala:27.28" *) 1'h0 : _001_;
  assign idMatch = & _007_;
  assign _092_ = & _091_;
  assign _079_ = & _078_;
  assign _047_ = & _046_;
  assign _015_ = & _014_;
  assign _019_ = & _018_;
  assign _085_ = & _084_;
  assign _069_ = & _068_;
  assign _074_ = & _073_;
  assign _057_ = & _056_;
  assign _067_ = & _066_;
  assign _026_ = & _025_;
  assign _035_ = & _034_;
  assign _041_ = & _040_;
  assign _005_ = _004_ ^ io_acceptanceCode_0;
  assign _089_ = _076_ ^ _087_;
  assign _094_ = io_data0 ^ io_acceptanceCode_2;
  assign _044_ = _076_ ^ _042_;
  assign _012_ = _050_ ^ io_acceptanceCode_2;
  assign _016_ = _070_ ^ io_acceptanceCode_3;
  assign _082_ = io_data1 ^ io_acceptanceCode_3;
  assign _051_ = _050_ ^ io_acceptanceCode_0;
  assign _071_ = _070_ ^ io_acceptanceCode_1;
  assign _054_ = _053_ ^ io_acceptanceCode_2;
  assign _064_ = _060_ ^ _061_;
  assign _023_ = _049_ ^ _021_;
  assign _032_ = _029_ ^ _030_;
  assign _038_ = _004_ ^ io_acceptanceCode_2;
  assign _004_ = io_id[10:3];
  assign _075_ = io_id[2:0];
  assign _076_ = { _075_, io_rtr1 };
  assign _087_ = io_acceptanceCode_1[7:4];
  assign _088_ = io_acceptanceMask_1[7:4];
  assign _050_ = io_id[28:21];
  assign _070_ = io_id[20:13];
  assign _053_ = io_id[12:5];
  assign _059_ = io_id[4:0];
  assign _060_ = { _059_, io_rtr2 };
  assign _061_ = io_acceptanceCode_3[7:2];
  assign _063_ = io_acceptanceMask_3[7:2];
  assign _049_ = io_data0[7:4];
  assign _021_ = io_acceptanceCode_1[3:0];
  assign _022_ = io_acceptanceMask_1[3:0];
  assign _029_ = io_data0[3:0];
  assign _030_ = io_acceptanceCode_3[3:0];
  assign _031_ = io_acceptanceMask_3[3:0];
  assign _042_ = io_acceptanceCode_3[7:4];
  assign _043_ = io_acceptanceMask_3[7:4];
  assign io_idOk = idOk;
  assign _096_ = reset;
  assign \idOk$process$CanAcf  = _095_;
endmodule

(* cells_not_processed =  1  *)
module CanBsp(clock, reset, io_samplePoint, io_sampledBit, io_sampledBitQ, io_txPoint, io_hardSync, io_addr, io_dataIn, io_dataOut, io_resetMode, io_listenOnlyMode, io_acceptanceFilterMode, io_extendedMode, io_selfTestMode, io_releaseBuffer, io_txRequest, io_abortTx, io_selfRxRequest, io_singleShotTransmission, io_txState
, io_txStateQ, io_overloadFrame, io_readArbitrationLostCaptureReg, io_readErrorCodeCaptureReg, io_errorCaptureCode, io_errorWarningLimit, io_writeEnReceiveErrorCounter, io_writeEnTransmitErrorCounter, io_rxIdle, io_transmitting, io_transmitter, io_goRxInter, io_notFirstBitOfInter, io_rxInter, io_setResetMode, io_nodeBusOff, io_errorStatus, io_rxErrorCount, io_txErrorCount, io_transmitStatus, io_receiveStatus
, io_txSuccessful, io_needToTx, io_overrun, io_infoEmpty, io_setBusErrorIrq, io_setArbitrationLostIrq, io_arbitrationLostCapture, io_nodeErrorPassive, io_nodeErrorActive, io_rxMessageCounter, io_acceptanceCode_0, io_acceptanceCode_1, io_acceptanceCode_2, io_acceptanceCode_3, io_acceptanceMask_0, io_acceptanceMask_1, io_acceptanceMask_2, io_acceptanceMask_3, io_txData_0, io_txData_1, io_txData_2
, io_txData_3, io_txData_4, io_txData_5, io_txData_6, io_txData_7, io_txData_8, io_txData_9, io_txData_10, io_txData_11, io_txData_12, io_tx, io_txNext, io_busOffOn, io_goOverloadFrame, io_goErrorFrame, io_goTx, io_sendAck);
  (* src = "CanBsp.scala:292.24|CanBsp.scala:293.12|CanBsp.scala:83.30" *)
  wire _0000_;
  (* src = "CanBsp.scala:290.35|CanBsp.scala:291.12" *)
  wire _0001_;
  (* src = "CanBsp.scala:322.24|CanBsp.scala:323.12|CanBsp.scala:116.30" *)
  wire _0002_;
  (* src = "CanBsp.scala:636.25|CanBsp.scala:637.21" *)
  wire _0003_;
  (* src = "CanBsp.scala:644.34|CanBsp.scala:645.19|CanBsp.scala:79.37" *)
  wire _0004_;
  (* src = "CanBsp.scala:642.46|CanBsp.scala:643.19" *)
  wire _0005_;
  (* src = "CanBsp.scala:650.67|CanBsp.scala:651.18|CanBsp.scala:151.36" *)
  wire [2:0] _0006_;
  (* src = "CanBsp.scala:648.67|CanBsp.scala:649.18" *)
  wire [2:0] _0007_;
  (* src = "CanBsp.scala:656.68|CanBsp.scala:657.24|CanBsp.scala:148.42" *)
  wire _0008_;
  (* src = "CanBsp.scala:654.67|CanBsp.scala:655.24" *)
  wire _0009_;
  (* src = "CanBsp.scala:662.46|CanBsp.scala:663.18|CanBsp.scala:152.36" *)
  wire [2:0] _0010_;
  (* src = "CanBsp.scala:660.67|CanBsp.scala:661.18" *)
  wire [2:0] _0011_;
  (* src = "CanBsp.scala:320.34|CanBsp.scala:321.12" *)
  wire _0012_;
  (* src = "CanBsp.scala:682.29|CanBsp.scala:690.19" *)
  wire _0013_;
  (* src = "CanBsp.scala:693.33|CanBsp.scala:694.19|CanBsp.scala:696.19" *)
  wire _0014_;
  (* src = "CanBsp.scala:701.30|CanBsp.scala:702.17|CanBsp.scala:704.17" *)
  wire _0015_;
  (* src = "CanBsp.scala:699.39|CanBsp.scala:700.19" *)
  wire _0016_;
  (* src = "CanBsp.scala:692.55" *)
  wire _0017_;
  (* src = "CanBsp.scala:681.41" *)
  wire _0018_;
  (* src = "CanBsp.scala:328.22|CanBsp.scala:329.10|CanBsp.scala:118.27" *)
  wire _0019_;
  (* src = "CanBsp.scala:710.26|CanBsp.scala:711.8|CanBsp.scala:103.26" *)
  wire _0020_;
  (* src = "CanBsp.scala:708.22|CanBsp.scala:709.8" *)
  wire _0021_;
  (* src = "CanBsp.scala:716.26|CanBsp.scala:717.9|CanBsp.scala:159.27" *)
  wire _0022_;
  (* src = "CanBsp.scala:714.22|CanBsp.scala:715.9" *)
  wire _0023_;
  (* src = "CanBsp.scala:725.27|CanBsp.scala:726.13|CanBsp.scala:728.13" *)
  wire _0024_;
  (* src = "CanBsp.scala:723.23|CanBsp.scala:724.13" *)
  wire _0025_;
  (* src = "CanBsp.scala:721.18|CanBsp.scala:722.13" *)
  wire _0026_;
  (* src = "CanBsp.scala:735.27|CanBsp.scala:736.13|CanBsp.scala:738.13" *)
  wire _0027_;
  (* src = "CanBsp.scala:733.23|CanBsp.scala:734.13" *)
  wire _0028_;
  (* src = "CanBsp.scala:326.34|CanBsp.scala:327.10" *)
  wire _0029_;
  (* src = "CanBsp.scala:731.18|CanBsp.scala:732.13" *)
  wire _0030_;
  (* src = "CanBsp.scala:744.81|CanBsp.scala:745.15|CanBsp.scala:164.33" *)
  wire [5:0] _0031_;
  (* src = "CanBsp.scala:742.22|CanBsp.scala:743.15" *)
  wire [5:0] _0032_;
  (* src = "CanBsp.scala:750.45|CanBsp.scala:751.14|CanBsp.scala:93.32" *)
  wire _0033_;
  (* src = "CanBsp.scala:748.130|CanBsp.scala:749.14" *)
  wire _0034_;
  (* src = "CanBsp.scala:758.25|CanBsp.scala:759.22|CanBsp.scala:126.40" *)
  wire _0035_;
  (* src = "CanBsp.scala:756.35|CanBsp.scala:757.22" *)
  wire _0036_;
  (* src = "CanBsp.scala:764.23|CanBsp.scala:765.13|CanBsp.scala:75.31" *)
  wire _0037_;
  (* src = "CanBsp.scala:762.68|CanBsp.scala:763.13" *)
  wire _0038_;
  (* src = "CanBsp.scala:334.22|CanBsp.scala:335.10|CanBsp.scala:117.28" *)
  wire _0039_;
  (* src = "CanBsp.scala:770.59|CanBsp.scala:771.17|CanBsp.scala:87.35" *)
  wire _0040_;
  (* src = "CanBsp.scala:768.17|CanBsp.scala:769.17" *)
  wire _0041_;
  (* src = "CanBsp.scala:776.98|CanBsp.scala:777.18|CanBsp.scala:85.36" *)
  wire _0042_;
  (* src = "CanBsp.scala:774.69|CanBsp.scala:775.18" *)
  wire _0043_;
  (* src = "CanBsp.scala:782.76|CanBsp.scala:783.13|CanBsp.scala:177.31" *)
  wire _0044_;
  (* src = "CanBsp.scala:780.63|CanBsp.scala:781.13" *)
  wire _0045_;
  (* src = "CanBsp.scala:788.57|CanBsp.scala:789.18|CanBsp.scala:178.36" *)
  wire _0046_;
  (* src = "CanBsp.scala:786.64|CanBsp.scala:787.18" *)
  wire _0047_;
  (* src = "CanBsp.scala:794.45|CanBsp.scala:795.16|CanBsp.scala:179.34" *)
  wire [2:0] _0048_;
  (* src = "CanBsp.scala:792.64|CanBsp.scala:793.16" *)
  wire [2:0] _0049_;
  (* src = "CanBsp.scala:332.35|CanBsp.scala:333.10" *)
  wire _0050_;
  (* src = "CanBsp.scala:800.26|CanBsp.scala:801.15|CanBsp.scala:166.33" *)
  wire _0051_;
  (* src = "CanBsp.scala:798.56|CanBsp.scala:799.15" *)
  wire _0052_;
  (* src = "CanBsp.scala:806.91|CanBsp.scala:807.21|CanBsp.scala:154.39" *)
  wire _0053_;
  (* src = "CanBsp.scala:804.36|CanBsp.scala:805.21" *)
  wire _0054_;
  (* src = "CanBsp.scala:810.24|CanBsp.scala:811.23|CanBsp.scala:156.41" *)
  wire _0055_;
  (* src = "CanBsp.scala:817.29|CanBsp.scala:818.22|CanBsp.scala:820.22" *)
  wire [4:0] _0056_;
  (* src = "CanBsp.scala:816.38|CanBsp.scala:157.38" *)
  wire [4:0] _0057_;
  (* src = "CanBsp.scala:824.34|CanBsp.scala:825.28|CanBsp.scala:99.46" *)
  wire [4:0] _0058_;
  (* src = "CanBsp.scala:830.40|CanBsp.scala:831.24|CanBsp.scala:158.42" *)
  wire _0059_;
  (* src = "CanBsp.scala:828.42|CanBsp.scala:829.24" *)
  wire _0060_;
  (* src = "CanBsp.scala:340.23|CanBsp.scala:341.11|CanBsp.scala:119.29" *)
  wire _0061_;
  (* src = "CanBsp.scala:841.39|CanBsp.scala:842.24|CanBsp.scala:844.24" *)
  wire [8:0] _0062_;
  (* src = "CanBsp.scala:850.116|CanBsp.scala:851.24|CanBsp.scala:95.36" *)
  wire [8:0] _0063_;
  (* src = "CanBsp.scala:847.40|CanBsp.scala:848.24" *)
  wire [8:0] _0064_;
  (* src = "CanBsp.scala:846.43|CanBsp.scala:95.36" *)
  wire [8:0] _0065_;
  (* src = "CanBsp.scala:840.83" *)
  wire [8:0] _0066_;
  (* src = "CanBsp.scala:839.68|CanBsp.scala:95.36" *)
  wire [8:0] _0067_;
  (* src = "CanBsp.scala:836.30|CanBsp.scala:837.18" *)
  wire [8:0] _0068_;
  (* src = "CanBsp.scala:834.58|CanBsp.scala:835.18" *)
  wire [8:0] _0069_;
  (* src = "CanBsp.scala:868.38|CanBsp.scala:869.22|CanBsp.scala:97.36" *)
  wire [8:0] _0070_;
  (* src = "CanBsp.scala:864.53|CanBsp.scala:97.36" *)
  wire [8:0] _0071_;
  (* src = "CanBsp.scala:338.46|CanBsp.scala:339.11" *)
  wire _0072_;
  (* src = "CanBsp.scala:862.68|CanBsp.scala:863.20" *)
  wire [8:0] _0073_;
  (* src = "CanBsp.scala:860.27|CanBsp.scala:861.20" *)
  wire [8:0] _0074_;
  (* src = "CanBsp.scala:857.40|CanBsp.scala:858.18" *)
  wire [8:0] _0075_;
  (* src = "CanBsp.scala:876.155|CanBsp.scala:877.22|CanBsp.scala:101.40" *)
  wire _0076_;
  (* src = "CanBsp.scala:874.57|CanBsp.scala:875.22" *)
  wire _0077_;
  (* src = "CanBsp.scala:884.101|CanBsp.scala:885.16|CanBsp.scala:91.34" *)
  wire _0078_;
  (* src = "CanBsp.scala:882.138|CanBsp.scala:883.16" *)
  wire _0079_;
  (* src = "CanBsp.scala:889.60|CanBsp.scala:890.18|CanBsp.scala:892.18" *)
  wire [3:0] _0080_;
  (* src = "CanBsp.scala:888.24|CanBsp.scala:167.34" *)
  wire [3:0] _0081_;
  (* src = "CanBsp.scala:898.87|CanBsp.scala:899.18|CanBsp.scala:168.36" *)
  wire _0082_;
  (* src = "CanBsp.scala:346.24|CanBsp.scala:347.12|CanBsp.scala:120.30" *)
  wire _0083_;
  (* src = "CanBsp.scala:896.68|CanBsp.scala:897.18" *)
  wire _0084_;
  (* src = "CanBsp.scala:910.43|CanBsp.scala:911.23|CanBsp.scala:169.41" *)
  wire _0085_;
  (* src = "CanBsp.scala:908.34|CanBsp.scala:909.23" *)
  wire _0086_;
  (* src = "CanBsp.scala:916.33|CanBsp.scala:917.22|CanBsp.scala:81.40" *)
  wire [7:0] _0087_;
  (* src = "CanBsp.scala:914.36|CanBsp.scala:915.22" *)
  wire [7:0] _0088_;
  (* src = "CanBsp.scala:929.24|CanBsp.scala:930.26|CanBsp.scala:932.26" *)
  wire [1:0] _0089_;
  (* src = "CanBsp.scala:927.23|CanBsp.scala:928.26" *)
  wire [1:0] _0090_;
  (* src = "CanBsp.scala:942.33|CanBsp.scala:943.29|CanBsp.scala:182.47" *)
  wire _0091_;
  (* src = "CanBsp.scala:344.35|CanBsp.scala:345.12" *)
  wire _0092_;
  (* src = "CanBsp.scala:940.36|CanBsp.scala:941.29" *)
  wire _0093_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0094_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0095_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0096_;
  (* src = "CanBsp.scala:244.63" *)
  wire [3:0] _0097_;
  (* src = "CanBsp.scala:244.37" *)
  wire [4:0] _0098_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0099_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0100_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0101_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0102_;
  (* src = "CanBsp.scala:298.23|CanBsp.scala:299.11|CanBsp.scala:112.29" *)
  wire _0103_;
  (* src = "CanBsp.scala:352.23|CanBsp.scala:353.11|CanBsp.scala:121.29" *)
  wire _0104_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0105_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0106_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0107_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0108_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0109_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0110_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0111_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0112_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0113_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0114_;
  (* src = "CanBsp.scala:350.38|CanBsp.scala:351.11" *)
  wire _0115_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0116_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0117_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0118_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0119_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0120_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0121_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0122_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0123_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0124_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0125_;
  (* src = "CanBsp.scala:358.26|CanBsp.scala:359.14|CanBsp.scala:122.32" *)
  wire _0126_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0127_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0128_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0129_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0130_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0131_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0132_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0133_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0134_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0135_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0136_;
  (* src = "CanBsp.scala:356.35|CanBsp.scala:357.14" *)
  wire _0137_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0138_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0139_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0140_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0141_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _0142_;
  (* src = "CanBsp.scala:946.58" *)
  wire [8:0] _0143_;
  (* src = "CanBsp.scala:160.31|CanBsp.scala:160.31" *)
  wire [4:0] _0144_;
  (* src = "CanBsp.scala:161.33|CanBsp.scala:161.33" *)
  wire [3:0] _0145_;
  (* src = "CanBsp.scala:364.23|CanBsp.scala:365.11|CanBsp.scala:123.29" *)
  wire _0146_;
  (* src = "CanBsp.scala:362.38|CanBsp.scala:363.11" *)
  wire _0147_;
  (* src = "CanBsp.scala:370.26|CanBsp.scala:371.14|CanBsp.scala:124.32" *)
  wire _0148_;
  (* src = "CanBsp.scala:368.35|CanBsp.scala:369.14" *)
  wire _0149_;
  (* src = "CanBsp.scala:376.23|CanBsp.scala:377.11|CanBsp.scala:125.29" *)
  wire _0150_;
  (* src = "CanBsp.scala:374.61|CanBsp.scala:375.11" *)
  wire _0151_;
  (* src = "CanBsp.scala:296.36|CanBsp.scala:297.11" *)
  wire _0152_;
  (* src = "CanBsp.scala:382.28|CanBsp.scala:383.13|CanBsp.scala:89.31" *)
  wire _0153_;
  (* src = "CanBsp.scala:380.67|CanBsp.scala:381.13" *)
  wire _0154_;
  (* src = "CanBsp.scala:386.56|CanBsp.scala:387.8|CanBsp.scala:108.26" *)
  wire [28:0] _0155_;
  (* src = "CanBsp.scala:390.47|CanBsp.scala:391.10|CanBsp.scala:127.28" *)
  wire _0156_;
  (* src = "CanBsp.scala:394.47|CanBsp.scala:395.10|CanBsp.scala:129.28" *)
  wire _0157_;
  (* src = "CanBsp.scala:398.46|CanBsp.scala:399.9|CanBsp.scala:128.27" *)
  wire _0158_;
  (* src = "CanBsp.scala:402.46|CanBsp.scala:403.13|CanBsp.scala:107.31" *)
  wire [3:0] _0159_;
  (* src = "CanBsp.scala:406.47|CanBsp.scala:407.13|CanBsp.scala:131.31" *)
  wire [7:0] _0160_;
  (* src = "CanBsp.scala:418.43|CanBsp.scala:419.13|CanBsp.scala:138.31" *)
  wire [2:0] _0161_;
  (* src = "CanBsp.scala:304.24|CanBsp.scala:305.12|CanBsp.scala:113.30" *)
  wire _0162_;
  (* src = "CanBsp.scala:416.28|CanBsp.scala:417.13" *)
  wire [2:0] _0163_;
  (* src = "CanBsp.scala:426.46|CanBsp.scala:427.11|CanBsp.scala:130.29" *)
  wire [14:0] _0164_;
  (* src = "CanBsp.scala:432.44|CanBsp.scala:433.12|CanBsp.scala:106.30" *)
  wire [5:0] _0165_;
  (* src = "CanBsp.scala:430.132|CanBsp.scala:431.12" *)
  wire [5:0] _0166_;
  (* src = "CanBsp.scala:438.23|CanBsp.scala:439.14|CanBsp.scala:141.30" *)
  wire [2:0] _0167_;
  (* src = "CanBsp.scala:302.35|CanBsp.scala:303.12" *)
  wire _0168_;
  (* src = "CanBsp.scala:436.63|CanBsp.scala:437.14" *)
  wire [2:0] _0169_;
  (* src = "CanBsp.scala:435.24|CanBsp.scala:141.30" *)
  wire [2:0] _0170_;
  (* src = "CanBsp.scala:445.31|CanBsp.scala:446.19|CanBsp.scala:139.37" *)
  wire _0171_;
  (* src = "CanBsp.scala:443.23|CanBsp.scala:444.19" *)
  wire _0172_;
  (* src = "CanBsp.scala:454.50|CanBsp.scala:455.19|CanBsp.scala:457.19" *)
  wire [2:0] _0173_;
  (* src = "CanBsp.scala:452.31|CanBsp.scala:453.19" *)
  wire [2:0] _0174_;
  (* src = "CanBsp.scala:451.46|CanBsp.scala:109.35" *)
  wire [2:0] _0175_;
  (* src = "CanBsp.scala:449.25|CanBsp.scala:450.17" *)
  wire [2:0] _0176_;
  (* src = "CanBsp.scala:466.31|CanBsp.scala:467.21|CanBsp.scala:469.21" *)
  wire [2:0] _0177_;
  (* src = "CanBsp.scala:464.33|CanBsp.scala:465.21" *)
  wire [2:0] _0178_;
  (* src = "CanBsp.scala:310.23|CanBsp.scala:311.11|CanBsp.scala:114.29" *)
  wire _0179_;
  (* src = "CanBsp.scala:463.40|CanBsp.scala:110.37" *)
  wire [2:0] _0180_;
  (* src = "CanBsp.scala:461.40|CanBsp.scala:462.19" *)
  wire [2:0] _0181_;
  (* src = "CanBsp.scala:475.27|CanBsp.scala:476.15|CanBsp.scala:140.33" *)
  wire _0182_;
  (* src = "CanBsp.scala:473.22|CanBsp.scala:474.15" *)
  wire _0183_;
  (* src = "CanBsp.scala:481.23|CanBsp.scala:482.12|CanBsp.scala:153.30" *)
  wire _0184_;
  (* src = "CanBsp.scala:479.40|CanBsp.scala:480.12" *)
  wire _0185_;
  (* src = "CanBsp.scala:487.22|CanBsp.scala:488.19|CanBsp.scala:172.37" *)
  wire _0186_;
  (* src = "CanBsp.scala:485.61|CanBsp.scala:486.19" *)
  wire _0187_;
  (* src = "CanBsp.scala:493.22|CanBsp.scala:494.19|CanBsp.scala:173.37" *)
  wire _0188_;
  (* src = "CanBsp.scala:491.61|CanBsp.scala:492.19" *)
  wire _0189_;
  (* src = "CanBsp.scala:308.45|CanBsp.scala:309.11" *)
  wire _0190_;
  (* src = "CanBsp.scala:499.84|CanBsp.scala:500.18|CanBsp.scala:176.38" *)
  wire _0191_;
  (* src = "CanBsp.scala:497.40|CanBsp.scala:498.18" *)
  wire _0192_;
  (* src = "CanBsp.scala:505.61|CanBsp.scala:506.18|CanBsp.scala:176.38" *)
  wire _0193_;
  (* src = "CanBsp.scala:503.38|CanBsp.scala:504.18" *)
  wire _0194_;
  (* src = "CanBsp.scala:511.24|CanBsp.scala:512.21|CanBsp.scala:174.39" *)
  wire _0195_;
  (* src = "CanBsp.scala:509.61|CanBsp.scala:510.21" *)
  wire _0196_;
  (* src = "CanBsp.scala:517.23|CanBsp.scala:518.20|CanBsp.scala:175.38" *)
  wire _0197_;
  (* src = "CanBsp.scala:515.61|CanBsp.scala:516.20" *)
  wire _0198_;
  (* src = "CanBsp.scala:547.89|CanBsp.scala:548.12|CanBsp.scala:162.30" *)
  wire _0199_;
  (* src = "CanBsp.scala:545.21|CanBsp.scala:546.12" *)
  wire _0200_;
  (* src = "CanBsp.scala:316.23|CanBsp.scala:317.11|CanBsp.scala:115.29" *)
  wire _0201_;
  (* src = "CanBsp.scala:553.38|CanBsp.scala:554.15|CanBsp.scala:161.33" *)
  wire [3:0] _0202_;
  (* src = "CanBsp.scala:551.21|CanBsp.scala:552.15" *)
  wire [3:0] _0203_;
  (* src = "CanBsp.scala:559.22|CanBsp.scala:560.13|CanBsp.scala:160.31" *)
  wire [4:0] _0204_;
  (* src = "CanBsp.scala:557.21|CanBsp.scala:558.13" *)
  wire [4:0] _0205_;
  (* src = "CanBsp.scala:592.31|CanBsp.scala:593.16|CanBsp.scala:143.34" *)
  wire _0206_;
  (* src = "CanBsp.scala:590.64|CanBsp.scala:591.16" *)
  wire _0207_;
  (* src = "CanBsp.scala:598.59|CanBsp.scala:599.15|CanBsp.scala:145.33" *)
  wire [2:0] _0208_;
  (* src = "CanBsp.scala:596.64|CanBsp.scala:597.15" *)
  wire [2:0] _0209_;
  (* src = "CanBsp.scala:604.29|CanBsp.scala:605.26|CanBsp.scala:180.44" *)
  wire _0210_;
  (* src = "CanBsp.scala:602.64|CanBsp.scala:603.26" *)
  wire _0211_;
  (* src = "CanBsp.scala:314.37|CanBsp.scala:315.11" *)
  wire _0212_;
  (* src = "CanBsp.scala:610.60|CanBsp.scala:611.21|CanBsp.scala:144.39" *)
  wire _0213_;
  (* src = "CanBsp.scala:608.64|CanBsp.scala:609.21" *)
  wire _0214_;
  (* src = "CanBsp.scala:616.44|CanBsp.scala:617.15|CanBsp.scala:146.33" *)
  wire [2:0] _0215_;
  (* src = "CanBsp.scala:614.64|CanBsp.scala:615.15" *)
  wire [2:0] _0216_;
  (* src = "CanBsp.scala:622.95|CanBsp.scala:623.24|CanBsp.scala:147.42" *)
  wire [2:0] _0217_;
  (* src = "CanBsp.scala:620.85|CanBsp.scala:621.24" *)
  wire [2:0] _0218_;
  (* src = "CanBsp.scala:629.78|CanBsp.scala:630.18|CanBsp.scala:632.18" *)
  wire [2:0] _0219_;
  (* src = "CanBsp.scala:628.51|CanBsp.scala:142.34" *)
  wire [2:0] _0220_;
  (* src = "CanBsp.scala:626.82|CanBsp.scala:627.16" *)
  wire [2:0] _0221_;
  (* src = "CanBsp.scala:638.30|CanBsp.scala:639.21|CanBsp.scala:183.39" *)
  wire _0222_;
  wire [2:0] _0223_;
  wire [7:0] _0224_;
  wire _0225_;
  wire [3:0] _0226_;
  wire [1:0] _0227_;
  wire [15:0] _0228_;
  wire [15:0] _0229_;
  wire [5:0] _0230_;
  wire [5:0] _0231_;
  wire [6:0] _0232_;
  wire [5:0] _0233_;
  wire [5:0] _0234_;
  wire [5:0] _0235_;
  wire [6:0] _0236_;
  wire [5:0] _0237_;
  wire [1:0] _0238_;
  wire [10:0] _0239_;
  wire [10:0] _0240_;
  wire [11:0] _0241_;
  wire [10:0] _0242_;
  wire [5:0] _0243_;
  wire [5:0] _0244_;
  wire [6:0] _0245_;
  wire [5:0] _0246_;
  wire [10:0] _0247_;
  wire [10:0] _0248_;
  wire [1:0] _0249_;
  wire [11:0] _0250_;
  wire [10:0] _0251_;
  wire [5:0] _0252_;
  wire [5:0] _0253_;
  wire [6:0] _0254_;
  wire [5:0] _0255_;
  wire [5:0] _0256_;
  wire [5:0] _0257_;
  wire [6:0] _0258_;
  wire [5:0] _0259_;
  wire [3:0] _0260_;
  wire [12:0] _0261_;
  wire [19:0] _0262_;
  wire [5:0] _0263_;
  wire [5:0] _0264_;
  wire [6:0] _0265_;
  wire [5:0] _0266_;
  wire [12:0] _0267_;
  wire [5:0] _0268_;
  wire [5:0] _0269_;
  wire [6:0] _0270_;
  wire [1:0] _0271_;
  wire [5:0] _0272_;
  wire [5:0] _0273_;
  wire [5:0] _0274_;
  wire [6:0] _0275_;
  wire [5:0] _0276_;
  wire [12:0] _0277_;
  wire [19:0] _0278_;
  wire [5:0] _0279_;
  wire [5:0] _0280_;
  wire [6:0] _0281_;
  wire [1:0] _0282_;
  wire [5:0] _0283_;
  wire [12:0] _0284_;
  wire [6:0] _0285_;
  wire [6:0] _0286_;
  wire [9:0] _0287_;
  wire [6:0] _0288_;
  wire [6:0] _0289_;
  wire [6:0] _0290_;
  wire [9:0] _0291_;
  wire [6:0] _0292_;
  wire [1:0] _0293_;
  wire [8:0] _0294_;
  wire [18:0] _0295_;
  wire [6:0] _0296_;
  wire [6:0] _0297_;
  wire [9:0] _0298_;
  wire [6:0] _0299_;
  wire [8:0] _0300_;
  wire [5:0] _0301_;
  wire [5:0] _0302_;
  wire [6:0] _0303_;
  wire [1:0] _0304_;
  wire [5:0] _0305_;
  wire [5:0] _0306_;
  wire [5:0] _0307_;
  wire [6:0] _0308_;
  wire [5:0] _0309_;
  wire [12:0] _0310_;
  wire [19:0] _0311_;
  wire [5:0] _0312_;
  wire [5:0] _0313_;
  wire [6:0] _0314_;
  wire [2:0] _0315_;
  wire [5:0] _0316_;
  wire [12:0] _0317_;
  wire [6:0] _0318_;
  wire [6:0] _0319_;
  wire [9:0] _0320_;
  wire [6:0] _0321_;
  wire [6:0] _0322_;
  wire [6:0] _0323_;
  wire [9:0] _0324_;
  wire [6:0] _0325_;
  wire [1:0] _0326_;
  wire [8:0] _0327_;
  wire [18:0] _0328_;
  wire [6:0] _0329_;
  wire [6:0] _0330_;
  wire [9:0] _0331_;
  wire [6:0] _0332_;
  wire [8:0] _0333_;
  wire [15:0] _0334_;
  wire [15:0] _0335_;
  wire [15:0] _0336_;
  wire [2:0] _0337_;
  wire [6:0] _0338_;
  wire [31:0] _0339_;
  wire [15:0] _0340_;
  wire [15:0] _0341_;
  wire [15:0] _0342_;
  wire [15:0] _0343_;
  wire [15:0] _0344_;
  wire [31:0] _0345_;
  wire [15:0] _0346_;
  wire [15:0] _0347_;
  wire [15:0] _0348_;
  wire [1:0] _0349_;
  wire [15:0] _0350_;
  wire [15:0] _0351_;
  wire [31:0] _0352_;
  wire [15:0] _0353_;
  wire [15:0] _0354_;
  wire [15:0] _0355_;
  wire [15:0] _0356_;
  wire [15:0] _0357_;
  wire [31:0] _0358_;
  wire [15:0] _0359_;
  wire [1:0] _0360_;
  wire [15:0] _0361_;
  wire [15:0] _0362_;
  wire [15:0] _0363_;
  wire [15:0] _0364_;
  wire [31:0] _0365_;
  wire [15:0] _0366_;
  wire [15:0] _0367_;
  wire [15:0] _0368_;
  wire [15:0] _0369_;
  wire [15:0] _0370_;
  wire [1:0] _0371_;
  wire [31:0] _0372_;
  wire [15:0] _0373_;
  wire [15:0] _0374_;
  wire [15:0] _0375_;
  wire [15:0] _0376_;
  wire [15:0] _0377_;
  wire [31:0] _0378_;
  wire [15:0] _0379_;
  wire [15:0] _0380_;
  wire [15:0] _0381_;
  wire [3:0] _0382_;
  wire [15:0] _0383_;
  wire [15:0] _0384_;
  wire [31:0] _0385_;
  wire [15:0] _0386_;
  wire [15:0] _0387_;
  wire [15:0] _0388_;
  wire [15:0] _0389_;
  wire [15:0] _0390_;
  wire [31:0] _0391_;
  wire [15:0] _0392_;
  wire [1:0] _0393_;
  wire [15:0] _0394_;
  wire [15:0] _0395_;
  wire [15:0] _0396_;
  wire [15:0] _0397_;
  wire [31:0] _0398_;
  wire [15:0] _0399_;
  wire [15:0] _0400_;
  wire [3:0] _0401_;
  wire [4:0] _0402_;
  wire [1:0] _0403_;
  wire [1:0] _0404_;
  wire [1:0] _0405_;
  wire [3:0] _0406_;
  wire [1:0] _0407_;
  wire [3:0] _0408_;
  wire [1:0] _0409_;
  wire [1:0] _0410_;
  wire [5:0] _0411_;
  wire [1:0] _0412_;
  wire [5:0] _0413_;
  wire [1:0] _0414_;
  wire [1:0] _0415_;
  wire [1:0] _0416_;
  wire [5:0] _0417_;
  wire [1:0] _0418_;
  wire [5:0] _0419_;
  wire [3:0] _0420_;
  wire [3:0] _0421_;
  wire [3:0] _0422_;
  wire [3:0] _0423_;
  wire [3:0] _0424_;
  wire [3:0] _0425_;
  wire [1:0] _0426_;
  wire [2:0] _0427_;
  wire [2:0] _0428_;
  wire [1:0] _0429_;
  wire [1:0] _0430_;
  wire [2:0] _0431_;
  wire [1:0] _0432_;
  wire [1:0] _0433_;
  wire [1:0] _0434_;
  wire [2:0] _0435_;
  wire [1:0] _0436_;
  wire [2:0] _0437_;
  wire [1:0] _0438_;
  wire [4:0] _0439_;
  wire [1:0] _0440_;
  wire [1:0] _0441_;
  wire [2:0] _0442_;
  wire [1:0] _0443_;
  wire [1:0] _0444_;
  wire [2:0] _0445_;
  wire [1:0] _0446_;
  wire [1:0] _0447_;
  wire _0448_;
  wire [1:0] _0449_;
  wire [2:0] _0450_;
  wire [1:0] _0451_;
  wire [1:0] _0452_;
  wire [1:0] _0453_;
  wire [2:0] _0454_;
  wire [1:0] _0455_;
  wire [1:0] _0456_;
  wire [4:0] _0457_;
  wire [1:0] _0458_;
  wire [1:0] _0459_;
  wire [1:0] _0460_;
  wire [2:0] _0461_;
  wire [1:0] _0462_;
  wire [1:0] _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire [5:0] _0469_;
  wire [1:0] _0470_;
  wire [1:0] _0471_;
  wire [3:0] _0472_;
  wire [1:0] _0473_;
  wire [1:0] _0474_;
  wire [1:0] _0475_;
  wire [1:0] _0476_;
  wire [1:0] _0477_;
  wire [1:0] _0478_;
  wire [3:0] _0479_;
  wire [1:0] _0480_;
  wire [1:0] _0481_;
  wire [1:0] _0482_;
  wire [1:0] _0483_;
  wire [2:0] _0484_;
  wire [1:0] _0485_;
  wire [6:0] _0486_;
  wire [1:0] _0487_;
  wire [1:0] _0488_;
  wire [1:0] _0489_;
  wire [1:0] _0490_;
  wire [3:0] _0491_;
  wire [1:0] _0492_;
  wire [1:0] _0493_;
  wire [1:0] _0494_;
  wire [1:0] _0495_;
  wire [2:0] _0496_;
  wire [1:0] _0497_;
  wire [5:0] _0498_;
  wire [5:0] _0499_;
  wire [1:0] _0500_;
  wire [9:0] _0501_;
  wire [5:0] _0502_;
  wire [5:0] _0503_;
  wire [5:0] _0504_;
  wire [9:0] _0505_;
  wire [5:0] _0506_;
  wire [8:0] _0507_;
  wire [5:0] _0508_;
  wire [5:0] _0509_;
  wire [9:0] _0510_;
  wire [3:0] _0511_;
  wire [5:0] _0512_;
  wire [8:0] _0513_;
  wire [15:0] _0514_;
  wire [15:0] _0515_;
  wire [15:0] _0516_;
  wire [31:0] _0517_;
  wire [15:0] _0518_;
  wire [15:0] _0519_;
  wire [15:0] _0520_;
  wire [15:0] _0521_;
  wire [1:0] _0522_;
  wire [15:0] _0523_;
  wire [31:0] _0524_;
  wire [15:0] _0525_;
  wire [15:0] _0526_;
  wire [15:0] _0527_;
  wire [15:0] _0528_;
  wire [15:0] _0529_;
  wire [31:0] _0530_;
  wire [15:0] _0531_;
  wire [15:0] _0532_;
  wire [1:0] _0533_;
  wire [15:0] _0534_;
  wire [15:0] _0535_;
  wire [15:0] _0536_;
  wire [31:0] _0537_;
  wire [15:0] _0538_;
  wire [15:0] _0539_;
  wire [15:0] _0540_;
  wire [15:0] _0541_;
  wire [15:0] _0542_;
  wire [31:0] _0543_;
  (* src = "CanBsp.scala:290.16" *)
  wire _0544_;
  (* src = "CanBsp.scala:296.17" *)
  wire _0545_;
  (* src = "CanBsp.scala:338.27" *)
  wire _0546_;
  (* src = "CanBsp.scala:598.38" *)
  wire _0547_;
  (* src = "CanBsp.scala:610.42" *)
  wire _0548_;
  (* src = "CanBsp.scala:610.25" *)
  wire _0549_;
  (* src = "CanBsp.scala:344.16" *)
  wire _0550_;
  (* src = "CanBsp.scala:616.30" *)
  wire _0551_;
  (* src = "CanBsp.scala:620.24" *)
  wire _0552_;
  (* src = "CanBsp.scala:620.42" *)
  wire _0553_;
  (* src = "CanBsp.scala:620.63" *)
  wire _0554_;
  (* src = "CanBsp.scala:622.68" *)
  wire _0555_;
  (* src = "CanBsp.scala:622.46" *)
  wire _0556_;
  (* src = "CanBsp.scala:350.19" *)
  wire _0557_;
  (* src = "CanBsp.scala:626.63" *)
  wire _0558_;
  (* src = "CanBsp.scala:628.43" *)
  wire _0559_;
  (* src = "CanBsp.scala:628.29" *)
  wire _0560_;
  (* src = "CanBsp.scala:629.21" *)
  wire _0561_;
  (* src = "CanBsp.scala:629.40" *)
  wire _0562_;
  (* src = "CanBsp.scala:642.27" *)
  wire _0563_;
  (* src = "CanBsp.scala:648.45" *)
  wire _0564_;
  (* src = "CanBsp.scala:650.31" *)
  wire _0565_;
  (* src = "CanBsp.scala:650.44" *)
  wire _0566_;
  (* src = "CanBsp.scala:656.51" *)
  wire _0567_;
  (* src = "CanBsp.scala:656.31" *)
  wire _0568_;
  (* src = "CanBsp.scala:362.19" *)
  wire _0569_;
  (* src = "CanBsp.scala:662.33" *)
  wire _0570_;
  (* src = "CanBsp.scala:678.22" *)
  wire _0571_;
  (* src = "CanBsp.scala:368.16" *)
  wire _0572_;
  (* src = "CanBsp.scala:682.22" *)
  wire _0573_;
  (* src = "CanBsp.scala:692.35" *)
  wire _0574_;
  (* src = "CanBsp.scala:693.26" *)
  wire _0575_;
  (* src = "CanBsp.scala:699.25" *)
  wire _0576_;
  (* src = "CanBsp.scala:744.52" *)
  wire _0577_;
  (* src = "CanBsp.scala:744.38" *)
  wire _0578_;
  (* src = "CanBsp.scala:744.63" *)
  wire _0579_;
  (* src = "CanBsp.scala:744.24" *)
  wire _0580_;
  (* src = "CanBsp.scala:748.24" *)
  wire _0581_;
  (* src = "CanBsp.scala:374.21" *)
  wire _0582_;
  (* src = "CanBsp.scala:748.53" *)
  wire _0583_;
  (* src = "CanBsp.scala:748.39" *)
  wire _0584_;
  (* src = "CanBsp.scala:748.87" *)
  wire _0585_;
  (* src = "CanBsp.scala:748.101" *)
  wire _0586_;
  (* src = "CanBsp.scala:748.73" *)
  wire _0587_;
  (* src = "CanBsp.scala:750.27" *)
  wire _0588_;
  (* src = "CanBsp.scala:756.21" *)
  wire _0589_;
  (* src = "CanBsp.scala:762.21" *)
  wire _0590_;
  (* src = "CanBsp.scala:374.39" *)
  wire _0591_;
  (* src = "CanBsp.scala:762.36" *)
  wire _0592_;
  (* src = "CanBsp.scala:762.49" *)
  wire _0593_;
  (* src = "CanBsp.scala:770.27" *)
  wire _0594_;
  (* src = "CanBsp.scala:770.48" *)
  wire _0595_;
  (* src = "CanBsp.scala:770.38" *)
  wire _0596_;
  (* src = "CanBsp.scala:774.24" *)
  wire _0597_;
  (* src = "CanBsp.scala:774.45" *)
  wire _0598_;
  (* src = "CanBsp.scala:774.55" *)
  wire _0599_;
  (* src = "CanBsp.scala:380.17" *)
  wire _0600_;
  (* src = "CanBsp.scala:776.49" *)
  wire _0601_;
  (* src = "CanBsp.scala:776.38" *)
  wire _0602_;
  (* src = "CanBsp.scala:776.83" *)
  wire _0603_;
  (* src = "CanBsp.scala:776.64" *)
  wire _0604_;
  (* src = "CanBsp.scala:780.21" *)
  wire _0605_;
  (* src = "CanBsp.scala:782.36" *)
  wire _0606_;
  (* src = "CanBsp.scala:782.53" *)
  wire _0607_;
  (* src = "CanBsp.scala:380.27" *)
  wire _0608_;
  (* src = "CanBsp.scala:788.22" *)
  wire _0609_;
  (* src = "CanBsp.scala:788.39" *)
  wire _0610_;
  (* src = "CanBsp.scala:794.27" *)
  wire _0611_;
  (* src = "CanBsp.scala:798.27" *)
  wire _0612_;
  (* src = "CanBsp.scala:302.16" *)
  wire _0613_;
  (* src = "CanBsp.scala:380.48" *)
  wire _0614_;
  (* src = "CanBsp.scala:798.40" *)
  wire _0615_;
  (* src = "CanBsp.scala:804.17" *)
  wire _0616_;
  (* src = "CanBsp.scala:806.29" *)
  wire _0617_;
  (* src = "CanBsp.scala:806.46" *)
  wire _0618_;
  (* src = "CanBsp.scala:806.54" *)
  wire _0619_;
  (* src = "CanBsp.scala:806.73" *)
  wire _0620_;
  (* src = "CanBsp.scala:386.32" *)
  wire _0621_;
  (* src = "CanBsp.scala:834.38" *)
  wire _0622_;
  (* src = "CanBsp.scala:839.48" *)
  wire _0623_;
  (* src = "CanBsp.scala:839.29" *)
  wire _0624_;
  (* src = "CanBsp.scala:840.23" *)
  wire _0625_;
  (* src = "CanBsp.scala:840.47" *)
  wire _0626_;
  (* src = "CanBsp.scala:840.44" *)
  wire _0627_;
  (* src = "CanBsp.scala:840.75" *)
  wire _0628_;
  (* src = "CanBsp.scala:386.23" *)
  wire _0629_;
  (* src = "CanBsp.scala:840.56" *)
  wire _0630_;
  (* src = "CanBsp.scala:841.30" *)
  wire _0631_;
  (* src = "CanBsp.scala:846.34" *)
  wire _0632_;
  (* src = "CanBsp.scala:847.32" *)
  wire _0633_;
  (* src = "CanBsp.scala:847.30" *)
  wire _0634_;
  (* src = "CanBsp.scala:849.38" *)
  wire _0635_;
  (* src = "CanBsp.scala:849.35" *)
  wire _0636_;
  (* src = "CanBsp.scala:849.61" *)
  wire _0637_;
  (* src = "CanBsp.scala:849.78" *)
  wire _0638_;
  (* src = "CanBsp.scala:849.97" *)
  wire _0639_;
  (* src = "CanBsp.scala:850.37" *)
  wire _0640_;
  (* src = "CanBsp.scala:849.119" *)
  wire _0641_;
  (* src = "CanBsp.scala:850.105" *)
  wire _0642_;
  (* src = "CanBsp.scala:850.83" *)
  wire _0643_;
  (* src = "CanBsp.scala:850.46" *)
  wire _0644_;
  (* src = "CanBsp.scala:862.30" *)
  wire _0645_;
  (* src = "CanBsp.scala:386.41" *)
  wire _0646_;
  (* src = "CanBsp.scala:862.56" *)
  wire _0647_;
  (* src = "CanBsp.scala:862.37" *)
  wire _0648_;
  (* src = "CanBsp.scala:864.31" *)
  wire _0649_;
  (* src = "CanBsp.scala:865.79" *)
  wire _0650_;
  (* src = "CanBsp.scala:390.23" *)
  wire _0651_;
  (* src = "CanBsp.scala:866.29" *)
  wire _0652_;
  (* src = "CanBsp.scala:866.26" *)
  wire _0653_;
  (* src = "CanBsp.scala:867.29" *)
  wire _0654_;
  (* src = "CanBsp.scala:867.40" *)
  wire _0655_;
  (* src = "CanBsp.scala:867.59" *)
  wire _0656_;
  (* src = "CanBsp.scala:867.76" *)
  wire _0657_;
  (* src = "CanBsp.scala:867.84" *)
  wire _0658_;
  (* src = "CanBsp.scala:867.12" *)
  wire _0659_;
  (* src = "CanBsp.scala:866.79" *)
  wire _0660_;
  (* src = "CanBsp.scala:865.107" *)
  wire _0661_;
  (* src = "CanBsp.scala:868.21" *)
  wire _0662_;
  (* src = "CanBsp.scala:867.106" *)
  wire _0663_;
  (* src = "CanBsp.scala:874.22" *)
  wire _0664_;
  (* src = "CanBsp.scala:874.47" *)
  wire _0665_;
  (* src = "CanBsp.scala:874.31" *)
  wire _0666_;
  (* src = "CanBsp.scala:876.29" *)
  wire _0667_;
  (* src = "CanBsp.scala:876.55" *)
  wire _0668_;
  (* src = "CanBsp.scala:390.32" *)
  wire _0669_;
  (* src = "CanBsp.scala:876.39" *)
  wire _0670_;
  (* src = "CanBsp.scala:876.121" *)
  wire _0671_;
  (* src = "CanBsp.scala:876.103" *)
  wire _0672_;
  (* src = "CanBsp.scala:876.66" *)
  wire _0673_;
  (* src = "CanBsp.scala:876.135" *)
  wire _0674_;
  (* src = "CanBsp.scala:882.25" *)
  wire _0675_;
  (* src = "CanBsp.scala:882.53" *)
  wire _0676_;
  (* src = "CanBsp.scala:394.23" *)
  wire _0677_;
  (* src = "CanBsp.scala:882.34" *)
  wire _0678_;
  (* src = "CanBsp.scala:882.62" *)
  wire _0679_;
  (* src = "CanBsp.scala:882.127" *)
  wire _0680_;
  (* src = "CanBsp.scala:882.114" *)
  wire _0681_;
  (* src = "CanBsp.scala:882.80" *)
  wire _0682_;
  (* src = "CanBsp.scala:884.31" *)
  wire _0683_;
  (* src = "CanBsp.scala:884.88" *)
  wire _0684_;
  (* src = "CanBsp.scala:884.75" *)
  wire _0685_;
  (* src = "CanBsp.scala:884.41" *)
  wire _0686_;
  (* src = "CanBsp.scala:889.24" *)
  wire _0687_;
  (* src = "CanBsp.scala:889.52" *)
  wire _0688_;
  (* src = "CanBsp.scala:889.39" *)
  wire _0689_;
  (* src = "CanBsp.scala:896.51" *)
  wire _0690_;
  (* src = "CanBsp.scala:896.37" *)
  wire _0691_;
  (* src = "CanBsp.scala:308.16" *)
  wire _0692_;
  (* src = "CanBsp.scala:394.32" *)
  wire _0693_;
  (* src = "CanBsp.scala:898.69" *)
  wire _0694_;
  (* src = "CanBsp.scala:398.23" *)
  wire _0695_;
  (* src = "CanBsp.scala:398.31" *)
  wire _0696_;
  (* src = "CanBsp.scala:402.23" *)
  wire _0697_;
  (* src = "CanBsp.scala:402.31" *)
  wire _0698_;
  (* src = "CanBsp.scala:406.23" *)
  wire _0699_;
  (* src = "CanBsp.scala:406.32" *)
  wire _0700_;
  (* src = "CanBsp.scala:308.26" *)
  wire _0701_;
  (* src = "CanBsp.scala:410.54" *)
  wire [2:0] _0702_;
  (* src = "CanBsp.scala:410.64" *)
  wire _0703_;
  (* src = "CanBsp.scala:410.46" *)
  wire _0704_;
  (* src = "CanBsp.scala:418.29" *)
  wire _0705_;
  (* src = "CanBsp.scala:426.23" *)
  wire _0706_;
  (* src = "CanBsp.scala:426.31" *)
  wire _0707_;
  (* src = "CanBsp.scala:314.18" *)
  wire _0708_;
  (* src = "CanBsp.scala:430.16" *)
  wire _0709_;
  (* src = "CanBsp.scala:430.26" *)
  wire _0710_;
  (* src = "CanBsp.scala:430.36" *)
  wire _0711_;
  (* src = "CanBsp.scala:430.47" *)
  wire _0712_;
  (* src = "CanBsp.scala:430.57" *)
  wire _0713_;
  (* src = "CanBsp.scala:430.67" *)
  wire _0714_;
  (* src = "CanBsp.scala:430.77" *)
  wire _0715_;
  (* src = "CanBsp.scala:430.92" *)
  wire _0716_;
  (* src = "CanBsp.scala:430.110" *)
  wire _0717_;
  (* src = "CanBsp.scala:320.15" *)
  wire _0718_;
  (* src = "CanBsp.scala:432.29" *)
  wire _0719_;
  (* src = "CanBsp.scala:461.21" *)
  wire _0720_;
  (* src = "CanBsp.scala:463.23" *)
  wire _0721_;
  (* src = "CanBsp.scala:466.22" *)
  wire _0722_;
  (* src = "CanBsp.scala:326.15" *)
  wire _0723_;
  (* src = "CanBsp.scala:479.21" *)
  wire _0724_;
  (* src = "CanBsp.scala:485.39" *)
  wire _0725_;
  (* src = "CanBsp.scala:497.24" *)
  wire _0726_;
  (* src = "CanBsp.scala:499.27" *)
  wire _0727_;
  (* src = "CanBsp.scala:499.47" *)
  wire _0728_;
  (* src = "CanBsp.scala:332.16" *)
  wire _0729_;
  (* src = "CanBsp.scala:499.64" *)
  wire _0730_;
  (* src = "CanBsp.scala:503.22" *)
  wire _0731_;
  (* src = "CanBsp.scala:505.29" *)
  wire _0732_;
  (* src = "CanBsp.scala:505.51" *)
  wire _0733_;
  (* src = "CanBsp.scala:547.27" *)
  wire _0734_;
  (* src = "CanBsp.scala:338.17" *)
  wire _0735_;
  (* src = "CanBsp.scala:547.34" *)
  wire _0736_;
  (* src = "CanBsp.scala:547.68" *)
  wire _0737_;
  (* src = "CanBsp.scala:547.53" *)
  wire _0738_;
  (* src = "CanBsp.scala:553.21" *)
  wire _0739_;
  (* src = "CanBsp.scala:590.24" *)
  wire _0740_;
  (* src = "CanBsp.scala:590.42" *)
  wire _0741_;
  (* src = "CanBsp.scala:596.24" *)
  wire _0742_;
  (* src = "CanBsp.scala:596.42" *)
  wire _0743_;
  (* src = "CanBsp.scala:598.25" *)
  wire _0744_;
  (* src = "CanBsp.scala:232.29" *)
  wire _0745_;
  (* src = "CanBsp.scala:232.46" *)
  wire _0746_;
  (* src = "CanBsp.scala:232.62" *)
  wire _0747_;
  (* src = "CanBsp.scala:232.78" *)
  wire _0748_;
  (* src = "CanBsp.scala:818.40" *)
  wire [5:0] _0749_;
  (* src = "CanBsp.scala:818.40" *)
  wire [4:0] _0750_;
  (* src = "CanBsp.scala:247.39" *)
  wire _0751_;
  (* src = "CanBsp.scala:247.48" *)
  wire _0752_;
  (* src = "CanBsp.scala:247.56" *)
  wire _0753_;
  (* src = "CanBsp.scala:253.41" *)
  wire [3:0] _0754_;
  (* src = "CanBsp.scala:253.68" *)
  wire [3:0] _0755_;
  (* src = "CanBsp.scala:433.22" *)
  wire [6:0] _0756_;
  (* src = "CanBsp.scala:433.22" *)
  wire [5:0] _0757_;
  (* src = "CanBsp.scala:215.40" *)
  wire _0758_;
  (* src = "CanBsp.scala:214.41" *)
  wire _0759_;
  (* src = "CanBsp.scala:225.66" *)
  wire [2:0] _0760_;
  (* src = "CanBsp.scala:225.71" *)
  wire [5:0] _0761_;
  (* src = "CanBsp.scala:225.85" *)
  wire [6:0] _0762_;
  (* src = "CanBsp.scala:225.85" *)
  wire [5:0] _0763_;
  (* src = "CanBsp.scala:261.38" *)
  wire _0764_;
  (* src = "CanBsp.scala:263.38" *)
  wire _0765_;
  (* src = "CanBsp.scala:263.73" *)
  wire _0766_;
  (* src = "CanBsp.scala:264.56" *)
  wire _0767_;
  (* src = "CanBsp.scala:264.39" *)
  wire _0768_;
  (* src = "CanBsp.scala:264.63" *)
  wire _0769_;
  (* src = "CanBsp.scala:264.60" *)
  wire _0770_;
  (* src = "CanBsp.scala:264.118" *)
  wire _0771_;
  (* src = "CanBsp.scala:264.102" *)
  wire _0772_;
  (* src = "CanBsp.scala:264.130" *)
  wire _0773_;
  (* src = "CanBsp.scala:264.127" *)
  wire _0774_;
  (* src = "CanBsp.scala:265.39" *)
  wire _0775_;
  (* src = "CanBsp.scala:265.81" *)
  wire _0776_;
  (* src = "CanBsp.scala:266.44" *)
  wire _0777_;
  (* src = "CanBsp.scala:269.25" *)
  wire _0778_;
  (* src = "CanBsp.scala:269.38" *)
  wire _0779_;
  (* src = "CanBsp.scala:269.146" *)
  wire _0780_;
  (* src = "CanBsp.scala:269.143" *)
  wire _0781_;
  (* src = "CanBsp.scala:269.162" *)
  wire _0782_;
  (* src = "CanBsp.scala:269.159" *)
  wire _0783_;
  (* src = "CanBsp.scala:269.178" *)
  wire _0784_;
  (* src = "CanBsp.scala:269.175" *)
  wire _0785_;
  (* src = "CanBsp.scala:269.194" *)
  wire _0786_;
  (* src = "CanBsp.scala:269.191" *)
  wire _0787_;
  (* src = "CanBsp.scala:269.210" *)
  wire _0788_;
  (* src = "CanBsp.scala:269.57" *)
  wire _0789_;
  (* src = "CanBsp.scala:269.66" *)
  wire _0790_;
  (* src = "CanBsp.scala:269.92" *)
  wire _0791_;
  (* src = "CanBsp.scala:269.83" *)
  wire _0792_;
  (* src = "CanBsp.scala:269.114" *)
  wire _0793_;
  (* src = "CanBsp.scala:269.111" *)
  wire _0794_;
  (* src = "CanBsp.scala:269.130" *)
  wire _0795_;
  (* src = "CanBsp.scala:269.127" *)
  wire _0796_;
  (* src = "CanBsp.scala:467.38" *)
  wire [3:0] _0797_;
  (* src = "CanBsp.scala:467.38" *)
  wire [2:0] _0798_;
  (* src = "CanBsp.scala:455.34" *)
  wire [3:0] _0799_;
  (* src = "CanBsp.scala:455.34" *)
  wire [2:0] _0800_;
  (* src = "CanBsp.scala:890.32" *)
  wire [4:0] _0801_;
  (* src = "CanBsp.scala:890.32" *)
  wire [3:0] _0802_;
  (* src = "CanBsp.scala:170.47" *)
  wire _0803_;
  (* src = "CanBsp.scala:170.77" *)
  wire _0804_;
  (* src = "CanBsp.scala:170.63" *)
  wire _0805_;
  (* src = "CanBsp.scala:170.87" *)
  wire _0806_;
  (* src = "CanBsp.scala:417.24" *)
  wire [3:0] _0807_;
  (* src = "CanBsp.scala:417.24" *)
  wire [2:0] _0808_;
  (* src = "CanBsp.scala:523.35" *)
  wire _0809_;
  (* src = "CanBsp.scala:482.21" *)
  wire _0810_;
  (* src = "CanBsp.scala:427.23" *)
  wire [13:0] _0811_;
  (* src = "Cat.scala:30.58" *)
  wire [14:0] _0812_;
  (* src = "CanBsp.scala:560.24" *)
  wire [4:0] _0813_;
  (* src = "Cat.scala:30.58" *)
  wire [3:0] _0814_;
  (* src = "CanBsp.scala:564.54" *)
  wire [4:0] _0815_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _0816_;
  (* src = "CanBsp.scala:571.28" *)
  wire [7:0] _0817_;
  (* src = "CanBsp.scala:572.32" *)
  wire [2:0] _0818_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _0819_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _0820_;
  (* src = "Lookup.scala:31.38" *)
  wire [5:0] _0821_;
  (* src = "Lookup.scala:31.38" *)
  wire _0822_;
  (* src = "CanBsp.scala:564.54" *)
  wire [3:0] _0823_;
  (* src = "Lookup.scala:31.38" *)
  wire _0824_;
  (* src = "Lookup.scala:31.38" *)
  wire _0825_;
  (* src = "Lookup.scala:31.38" *)
  wire _0826_;
  (* src = "Lookup.scala:31.38" *)
  wire _0827_;
  (* src = "Lookup.scala:31.38" *)
  wire _0828_;
  (* src = "Lookup.scala:31.38" *)
  wire _0829_;
  (* src = "Lookup.scala:31.38" *)
  wire _0830_;
  (* src = "Lookup.scala:31.38" *)
  wire _0831_;
  (* src = "Lookup.scala:31.38" *)
  wire _0832_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0833_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0834_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0835_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _0836_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0837_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0838_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0839_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0840_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0841_;
  (* src = "Lookup.scala:33.37" *)
  wire [7:0] _0842_;
  (* src = "CanBsp.scala:566.28" *)
  wire [7:0] _0843_;
  (* src = "CanBsp.scala:567.28" *)
  wire [7:0] _0844_;
  (* src = "CanBsp.scala:568.28" *)
  wire [7:0] _0845_;
  (* src = "CanBsp.scala:569.32" *)
  wire [4:0] _0846_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _0847_;
  (* src = "Cat.scala:30.58" *)
  wire [3:0] _0848_;
  (* src = "CanBsp.scala:623.46" *)
  wire [3:0] _0849_;
  (* src = "CanBsp.scala:623.46" *)
  wire [2:0] _0850_;
  (* src = "CanBsp.scala:439.24" *)
  wire [3:0] _0851_;
  (* src = "CanBsp.scala:439.24" *)
  wire [2:0] _0852_;
  (* src = "CanBsp.scala:245.28" *)
  wire _0853_;
  (* src = "CanBsp.scala:245.39" *)
  wire _0854_;
  (* src = "CanBsp.scala:245.48" *)
  wire _0855_;
  (* src = "CanBsp.scala:245.57" *)
  wire _0856_;
  (* src = "CanBsp.scala:245.74" *)
  wire _0857_;
  (* src = "CanBsp.scala:245.92" *)
  wire _0858_;
  (* src = "CanBsp.scala:245.108" *)
  wire _0859_;
  (* src = "CanBsp.scala:919.43" *)
  wire _0860_;
  (* src = "CanBsp.scala:919.51" *)
  wire _0861_;
  (* src = "CanBsp.scala:920.46" *)
  wire _0862_;
  (* src = "CanBsp.scala:920.53" *)
  wire _0863_;
  (* src = "CanBsp.scala:920.61" *)
  wire _0864_;
  (* src = "CanBsp.scala:920.70" *)
  wire _0865_;
  (* src = "CanBsp.scala:920.78" *)
  wire _0866_;
  (* src = "CanBsp.scala:920.89" *)
  wire _0867_;
  (* src = "CanBsp.scala:920.97" *)
  wire _0868_;
  (* src = "CanBsp.scala:920.108" *)
  wire _0869_;
  (* src = "CanBsp.scala:920.116" *)
  wire _0870_;
  (* src = "CanBsp.scala:921.22" *)
  wire _0871_;
  (* src = "CanBsp.scala:919.62" *)
  wire _0872_;
  (* src = "CanBsp.scala:921.12" *)
  wire _0873_;
  (* src = "CanBsp.scala:921.30" *)
  wire _0874_;
  (* src = "CanBsp.scala:921.39" *)
  wire _0875_;
  (* src = "CanBsp.scala:921.47" *)
  wire _0876_;
  (* src = "CanBsp.scala:921.55" *)
  wire _0877_;
  (* src = "CanBsp.scala:921.64" *)
  wire _0878_;
  (* src = "CanBsp.scala:921.71" *)
  wire _0879_;
  (* src = "CanBsp.scala:921.106" *)
  wire _0880_;
  (* src = "CanBsp.scala:922.13" *)
  wire _0881_;
  (* src = "CanBsp.scala:919.70" *)
  wire _0882_;
  (* src = "CanBsp.scala:922.21" *)
  wire _0883_;
  (* src = "CanBsp.scala:922.29" *)
  wire _0884_;
  (* src = "CanBsp.scala:922.37" *)
  wire _0885_;
  (* src = "CanBsp.scala:922.46" *)
  wire _0886_;
  (* src = "CanBsp.scala:922.57" *)
  wire _0887_;
  (* src = "CanBsp.scala:922.65" *)
  wire _0888_;
  (* src = "CanBsp.scala:922.78" *)
  wire _0889_;
  (* src = "CanBsp.scala:923.15" *)
  wire _0890_;
  (* src = "CanBsp.scala:923.42" *)
  wire _0891_;
  (* src = "CanBsp.scala:919.83" *)
  wire _0892_;
  (* src = "CanBsp.scala:923.32" *)
  wire _0893_;
  (* src = "CanBsp.scala:923.23" *)
  wire _0894_;
  (* src = "CanBsp.scala:923.51" *)
  wire _0895_;
  (* src = "CanBsp.scala:923.58" *)
  wire _0896_;
  (* src = "CanBsp.scala:923.65" *)
  wire _0897_;
  (* src = "CanBsp.scala:923.73" *)
  wire _0898_;
  (* src = "CanBsp.scala:923.81" *)
  wire _0899_;
  (* src = "CanBsp.scala:923.105" *)
  wire _0900_;
  (* src = "CanBsp.scala:923.92" *)
  wire _0901_;
  (* src = "CanBsp.scala:919.96" *)
  wire _0902_;
  (* src = "CanBsp.scala:920.22" *)
  wire _0903_;
  (* src = "CanBsp.scala:920.12" *)
  wire _0904_;
  (* src = "CanBsp.scala:920.30" *)
  wire _0905_;
  (* src = "CanBsp.scala:920.39" *)
  wire _0906_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _0907_;
  (* src = "CanBsp.scala:599.28" *)
  wire [3:0] _0908_;
  (* src = "CanBsp.scala:599.28" *)
  wire [2:0] _0909_;
  (* src = "CanBsp.scala:617.28" *)
  wire [3:0] _0910_;
  (* src = "CanBsp.scala:617.28" *)
  wire [2:0] _0911_;
  (* src = "CanBsp.scala:267.32" *)
  wire _0912_;
  (* src = "CanBsp.scala:267.54" *)
  wire _0913_;
  (* src = "CanBsp.scala:267.71" *)
  wire _0914_;
  (* src = "CanBsp.scala:267.114" *)
  wire _0915_;
  (* src = "CanBsp.scala:267.145" *)
  wire _0916_;
  (* src = "CanBsp.scala:267.131" *)
  wire _0917_;
  (* src = "CanBsp.scala:267.92" *)
  wire _0918_;
  (* src = "CanBsp.scala:229.47" *)
  wire _0919_;
  (* src = "CanBsp.scala:256.89" *)
  wire [4:0] _0920_;
  (* src = "CanBsp.scala:256.123" *)
  wire [4:0] _0921_;
  (* src = "CanBsp.scala:255.47" *)
  wire [3:0] _0922_;
  (* src = "CanBsp.scala:255.74" *)
  wire _0923_;
  (* src = "CanBsp.scala:255.89" *)
  wire [2:0] _0924_;
  (* src = "CanBsp.scala:222.57" *)
  wire _0925_;
  (* src = "CanBsp.scala:223.60" *)
  wire _0926_;
  (* src = "CanBsp.scala:223.82" *)
  wire _0927_;
  (* src = "CanBsp.scala:223.79" *)
  wire _0928_;
  (* src = "CanBsp.scala:223.35" *)
  wire _0929_;
  (* src = "CanBsp.scala:223.109" *)
  wire _0930_;
  (* src = "CanBsp.scala:223.128" *)
  wire _0931_;
  (* src = "CanBsp.scala:223.100" *)
  wire _0932_;
  (* src = "CanBsp.scala:222.68" *)
  wire _0933_;
  (* src = "CanBsp.scala:223.15" *)
  wire _0934_;
  (* src = "CanBsp.scala:222.88" *)
  wire _0935_;
  (* src = "CanBsp.scala:223.46" *)
  wire _0936_;
  (* src = "CanBsp.scala:223.52" *)
  wire _0937_;
  (* src = "CanBsp.scala:217.27" *)
  wire _0938_;
  (* src = "CanBsp.scala:217.47" *)
  wire _0939_;
  (* src = "CanBsp.scala:217.130" *)
  wire _0940_;
  (* src = "CanBsp.scala:217.64" *)
  wire _0941_;
  (* src = "CanBsp.scala:217.61" *)
  wire _0942_;
  (* src = "CanBsp.scala:217.80" *)
  wire _0943_;
  (* src = "CanBsp.scala:217.103" *)
  wire _0944_;
  (* src = "CanBsp.scala:217.89" *)
  wire _0945_;
  (* src = "CanBsp.scala:217.77" *)
  wire _0946_;
  (* src = "CanBsp.scala:217.113" *)
  wire _0947_;
  (* src = "CanBsp.scala:205.58" *)
  wire _0948_;
  (* src = "CanBsp.scala:205.81" *)
  wire _0949_;
  (* src = "CanBsp.scala:227.122" *)
  wire _0950_;
  (* src = "CanBsp.scala:227.78" *)
  wire _0951_;
  (* src = "CanBsp.scala:227.143" *)
  wire _0952_;
  (* src = "CanBsp.scala:227.134" *)
  wire _0953_;
  (* src = "CanBsp.scala:227.54" *)
  wire _0954_;
  (* src = "CanBsp.scala:227.101" *)
  wire _0955_;
  (* src = "CanBsp.scala:227.98" *)
  wire _0956_;
  (* src = "CanBsp.scala:226.120" *)
  wire _0957_;
  (* src = "CanBsp.scala:226.46" *)
  wire _0958_;
  (* src = "CanBsp.scala:226.69" *)
  wire _0959_;
  (* src = "CanBsp.scala:226.54" *)
  wire _0960_;
  (* src = "CanBsp.scala:226.104" *)
  wire [2:0] _0961_;
  (* src = "CanBsp.scala:226.113" *)
  wire _0962_;
  (* src = "CanBsp.scala:226.95" *)
  wire _0963_;
  (* src = "CanBsp.scala:226.78" *)
  wire _0964_;
  (* src = "CanBsp.scala:195.41" *)
  wire _0965_;
  (* src = "CanBsp.scala:195.39" *)
  wire _0966_;
  (* src = "CanBsp.scala:195.69" *)
  wire _0967_;
  (* src = "CanBsp.scala:198.55" *)
  wire _0968_;
  (* src = "CanBsp.scala:194.56" *)
  wire _0969_;
  (* src = "CanBsp.scala:194.85" *)
  wire _0970_;
  (* src = "CanBsp.scala:194.83" *)
  wire _0971_;
  (* src = "CanBsp.scala:201.63" *)
  wire _0972_;
  (* src = "CanBsp.scala:201.82" *)
  wire _0973_;
  (* src = "CanBsp.scala:196.26" *)
  wire _0974_;
  (* src = "CanBsp.scala:196.39" *)
  wire _0975_;
  (* src = "CanBsp.scala:196.56" *)
  wire _0976_;
  (* src = "CanBsp.scala:196.73" *)
  wire [3:0] _0977_;
  (* src = "CanBsp.scala:196.79" *)
  wire _0978_;
  (* src = "CanBsp.scala:199.56" *)
  wire _0979_;
  (* src = "CanBsp.scala:199.73" *)
  wire [4:0] _0980_;
  (* src = "CanBsp.scala:199.79" *)
  wire _0981_;
  (* src = "CanBsp.scala:554.28" *)
  wire [3:0] _0982_;
  (* src = "CanBsp.scala:241.50" *)
  wire [2:0] _0983_;
  (* src = "CanBsp.scala:387.17" *)
  wire [27:0] _0984_;
  (* src = "Cat.scala:30.58" *)
  wire [28:0] _0985_;
  (* src = "CanBsp.scala:946.58" *)
  wire _0986_;
  (* src = "CanBsp.scala:946.102" *)
  wire _0987_;
  (* src = "CanBsp.scala:946.83" *)
  wire _0988_;
  (* src = "CanBsp.scala:947.58" *)
  wire _0989_;
  (* src = "CanBsp.scala:947.86" *)
  wire _0990_;
  (* src = "CanBsp.scala:947.67" *)
  wire _0991_;
  (* src = "CanBsp.scala:286.70" *)
  wire _0992_;
  (* src = "CanBsp.scala:283.60" *)
  wire _0993_;
  (* src = "CanBsp.scala:283.88" *)
  wire _0994_;
  (* src = "CanBsp.scala:283.73" *)
  wire _0995_;
  (* src = "CanBsp.scala:282.171" *)
  wire _0996_;
  (* src = "CanBsp.scala:284.82" *)
  wire _0997_;
  (* src = "CanBsp.scala:284.60" *)
  wire _0998_;
  (* src = "CanBsp.scala:282.92" *)
  wire _0999_;
  (* src = "CanBsp.scala:282.112" *)
  wire _1000_;
  (* src = "CanBsp.scala:282.131" *)
  wire _1001_;
  (* src = "CanBsp.scala:282.149" *)
  wire _1002_;
  (* src = "CanBsp.scala:282.83" *)
  wire _1003_;
  (* src = "CanBsp.scala:235.36" *)
  wire _1004_;
  (* src = "CanBsp.scala:235.56" *)
  wire _1005_;
  (* src = "CanBsp.scala:235.46" *)
  wire _1006_;
  (* src = "CanBsp.scala:235.66" *)
  wire _1007_;
  (* src = "CanBsp.scala:754.95" *)
  wire _1008_;
  (* src = "CanBsp.scala:754.77" *)
  wire _1009_;
  (* src = "CanBsp.scala:754.65" *)
  wire _1010_;
  (* src = "CanBsp.scala:754.133" *)
  wire _1011_;
  (* src = "CanBsp.scala:880.47" *)
  wire _1012_;
  (* src = "CanBsp.scala:285.57" *)
  wire _1013_;
  (* src = "CanBsp.scala:936.67" *)
  wire _1014_;
  (* src = "CanBsp.scala:936.79" *)
  wire _1015_;
  (* src = "CanBsp.scala:936.63" *)
  wire _1016_;
  (* src = "CanBsp.scala:937.46" *)
  wire _1017_;
  (* src = "CanBsp.scala:937.66" *)
  wire _1018_;
  (* src = "CanBsp.scala:937.82" *)
  wire _1019_;
  (* src = "CanBsp.scala:260.31" *)
  wire _1020_;
  (* src = "CanBsp.scala:260.42" *)
  wire _1021_;
  (* src = "CanBsp.scala:260.39" *)
  wire _1022_;
  (* src = "CanBsp.scala:814.48" *)
  wire _1023_;
  (* src = "CanBsp.scala:814.45" *)
  wire _1024_;
  (* src = "CanBsp.scala:814.69" *)
  wire _1025_;
  (* src = "CanBsp.scala:938.43" *)
  wire _1026_;
  (* src = "CanBsp.scala:287.35" *)
  wire _1027_;
  (* src = "CanBsp.scala:935.60" *)
  wire _1028_;
  (* src = "CanBsp.scala:700.39" *)
  wire _1029_;
  (* src = "CanBsp.scala:700.67" *)
  wire _1030_;
  (* src = "CanBsp.scala:700.64" *)
  wire _1031_;
  (* src = "CanBsp.scala:700.48" *)
  wire _1032_;
  (* src = "CanBsp.scala:288.34" *)
  wire _1033_;
  (* src = "CanBsp.scala:288.49" *)
  wire _1034_;
  (* src = "CanBsp.scala:288.73" *)
  wire _1035_;
  (* src = "CanBsp.scala:288.70" *)
  wire _1036_;
  (* src = "CanBsp.scala:288.94" *)
  wire _1037_;
  (* src = "CanBsp.scala:288.91" *)
  wire _1038_;
  (* src = "CanBsp.scala:288.118" *)
  wire _1039_;
  (* src = "CanBsp.scala:192.48" *)
  wire [1:0] _1040_;
  (* src = "CanBsp.scala:192.54" *)
  wire _1041_;
  (* src = "CanBsp.scala:243.85" *)
  wire [4:0] _1042_;
  (* src = "CanBsp.scala:243.85" *)
  wire [3:0] _1043_;
  (* src = "CanBsp.scala:243.61" *)
  wire [3:0] _1044_;
  (* src = "CanBsp.scala:221.43" *)
  wire _1045_;
  (* src = "CanBsp.scala:271.48" *)
  wire _1046_;
  (* src = "CanBsp.scala:271.74" *)
  wire [2:0] _1047_;
  (* src = "CanBsp.scala:271.80" *)
  wire [5:0] _1048_;
  (* src = "CanBsp.scala:271.95" *)
  wire [6:0] _1049_;
  (* src = "CanBsp.scala:271.95" *)
  wire [5:0] _1050_;
  (* src = "CanBsp.scala:272.48" *)
  wire _1051_;
  (* src = "CanBsp.scala:272.74" *)
  wire [2:0] _1052_;
  (* src = "CanBsp.scala:272.80" *)
  wire [5:0] _1053_;
  (* src = "CanBsp.scala:272.95" *)
  wire [6:0] _1054_;
  (* src = "CanBsp.scala:272.95" *)
  wire [5:0] _1055_;
  (* src = "CanBsp.scala:238.40" *)
  wire _1056_;
  (* src = "CanBsp.scala:239.40" *)
  wire _1057_;
  (* src = "CanBsp.scala:651.34" *)
  wire [3:0] _1058_;
  (* src = "CanBsp.scala:651.34" *)
  wire [2:0] _1059_;
  (* src = "CanBsp.scala:663.34" *)
  wire [3:0] _1060_;
  (* src = "CanBsp.scala:663.34" *)
  wire [2:0] _1061_;
  (* src = "CanBsp.scala:268.48" *)
  wire _1062_;
  (* src = "CanBsp.scala:230.49" *)
  wire _1063_;
  (* src = "CanBsp.scala:630.32" *)
  wire [3:0] _1064_;
  (* src = "CanBsp.scala:630.32" *)
  wire [2:0] _1065_;
  (* src = "Bitwise.scala:109.18" *)
  wire [7:0] _1066_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1067_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1068_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1069_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1070_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1071_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1072_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1073_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1074_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1075_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1076_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1077_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1078_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1079_;
  (* src = "Bitwise.scala:109.44" *)
  wire [6:0] _1080_;
  (* src = "Bitwise.scala:109.18" *)
  wire [3:0] _1081_;
  (* src = "Bitwise.scala:109.18" *)
  wire [1:0] _1082_;
  (* src = "Bitwise.scala:109.18" *)
  wire _1083_;
  (* src = "Bitwise.scala:109.44" *)
  wire _1084_;
  (* src = "Bitwise.scala:109.44" *)
  wire [1:0] _1085_;
  (* src = "Bitwise.scala:109.18" *)
  wire _1086_;
  (* src = "Bitwise.scala:109.44" *)
  wire _1087_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1088_;
  (* src = "Bitwise.scala:109.44" *)
  wire [2:0] _1089_;
  (* src = "Bitwise.scala:109.18" *)
  wire [1:0] _1090_;
  (* src = "Bitwise.scala:109.18" *)
  wire _1091_;
  (* src = "Bitwise.scala:109.44" *)
  wire _1092_;
  (* src = "Bitwise.scala:109.44" *)
  wire _1093_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1094_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1095_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1096_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1097_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1098_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1099_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1100_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1101_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1102_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1103_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1104_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1105_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1106_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1107_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1108_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1109_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1110_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1111_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1112_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1113_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1114_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1115_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1116_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1117_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1118_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1119_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1120_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1121_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1122_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1123_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1124_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1125_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1126_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1127_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1128_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1129_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1130_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1131_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1132_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1133_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1134_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1135_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1136_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1137_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1138_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1139_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1140_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1141_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1142_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1143_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1144_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1145_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1146_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1147_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1148_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1149_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1150_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1151_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1152_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1153_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1154_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1155_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1156_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1157_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1158_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1159_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1160_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1161_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1162_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1163_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1164_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1165_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1166_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1167_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1168_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1169_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1170_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1171_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1172_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1173_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1174_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1175_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1176_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1177_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1178_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1179_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1180_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1181_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1182_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1183_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1184_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1185_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1186_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1187_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1188_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1189_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1190_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1191_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1192_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1193_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1194_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1195_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1196_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1197_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1198_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1199_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1200_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1201_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1202_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1203_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1204_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1205_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1206_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1207_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1208_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1209_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1210_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1211_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1212_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1213_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1214_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1215_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1216_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1217_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1218_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1219_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1220_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1221_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1222_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1223_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1224_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1225_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1226_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1227_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1228_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1229_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1230_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1231_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1232_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1233_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1234_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1235_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1236_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1237_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1238_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1239_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1240_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1241_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1242_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1243_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1244_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1245_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1246_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1247_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1248_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1249_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1250_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1251_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1252_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1253_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1254_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1255_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1256_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1257_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1258_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1259_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1260_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1261_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1262_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1263_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1264_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1265_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1266_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1267_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1268_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1269_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1270_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1271_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1272_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1273_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1274_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1275_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1276_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1277_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1278_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1279_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1280_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1281_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1282_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1283_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1284_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1285_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1286_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1287_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1288_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1289_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1290_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1291_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1292_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1293_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1294_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1295_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1296_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1297_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1298_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1299_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1300_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1301_;
  (* src = "Bitwise.scala:103.46" *)
  wire [5:0] _1302_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1303_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1304_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1305_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1306_;
  (* src = "Bitwise.scala:103.21" *)
  wire [6:0] _1307_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1308_;
  (* src = "Bitwise.scala:103.46" *)
  wire [6:0] _1309_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1310_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1311_;
  (* src = "Bitwise.scala:103.21" *)
  wire [3:0] _1312_;
  (* src = "Bitwise.scala:103.31" *)
  wire [7:0] _1313_;
  (* src = "Bitwise.scala:103.46" *)
  wire [3:0] _1314_;
  (* src = "Bitwise.scala:103.65" *)
  wire [7:0] _1315_;
  (* src = "Bitwise.scala:103.75" *)
  wire [7:0] _1316_;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] _1317_;
  (* src = "Bitwise.scala:103.21" *)
  wire [5:0] _1318_;
  (* src = "CanBsp.scala:209.27" *)
  wire _1319_;
  (* src = "CanBsp.scala:209.33" *)
  wire _1320_;
  (* src = "CanBsp.scala:209.48" *)
  wire _1321_;
  (* src = "CanBsp.scala:244.63" *)
  wire [4:0] _1322_;
  (* src = "CanBsp.scala:244.37" *)
  wire _1323_;
  (* src = "CanBsp.scala:274.31" *)
  wire _1324_;
  (* src = "CanBsp.scala:274.46" *)
  wire _1325_;
  (* src = "CanBsp.scala:275.93" *)
  wire _1326_;
  (* src = "CanBsp.scala:275.91" *)
  wire _1327_;
  (* src = "CanBsp.scala:275.120" *)
  wire _1328_;
  (* src = "CanBsp.scala:275.108" *)
  wire _1329_;
  (* src = "CanBsp.scala:274.130" *)
  wire _1330_;
  (* src = "CanBsp.scala:274.62" *)
  wire _1331_;
  (* src = "CanBsp.scala:276.74" *)
  wire _1332_;
  (* src = "CanBsp.scala:276.71" *)
  wire _1333_;
  (* src = "CanBsp.scala:276.106" *)
  wire _1334_;
  (* src = "CanBsp.scala:275.130" *)
  wire _1335_;
  (* src = "CanBsp.scala:274.59" *)
  wire _1336_;
  (* src = "CanBsp.scala:277.59" *)
  wire _1337_;
  (* src = "CanBsp.scala:277.71" *)
  wire _1338_;
  (* src = "CanBsp.scala:277.118" *)
  wire _1339_;
  (* src = "CanBsp.scala:277.106" *)
  wire _1340_;
  (* src = "CanBsp.scala:276.128" *)
  wire _1341_;
  (* src = "CanBsp.scala:274.71" *)
  wire _1342_;
  (* src = "CanBsp.scala:278.71" *)
  wire _1343_;
  (* src = "CanBsp.scala:278.118" *)
  wire _1344_;
  (* src = "CanBsp.scala:278.106" *)
  wire _1345_;
  (* src = "CanBsp.scala:277.139" *)
  wire _1346_;
  (* src = "CanBsp.scala:279.59" *)
  wire _1347_;
  (* src = "CanBsp.scala:278.139" *)
  wire _1348_;
  (* src = "CanBsp.scala:280.39" *)
  wire _1349_;
  (* src = "CanBsp.scala:280.52" *)
  wire _1350_;
  (* src = "CanBsp.scala:280.67" *)
  wire _1351_;
  (* src = "CanBsp.scala:274.104" *)
  wire _1352_;
  (* src = "CanBsp.scala:274.91" *)
  wire _1353_;
  (* src = "CanBsp.scala:274.120" *)
  wire _1354_;
  (* src = "CanBsp.scala:274.108" *)
  wire _1355_;
  (* src = "CanBsp.scala:270.49" *)
  wire _1356_;
  (* src = "CanBsp.scala:270.62" *)
  wire _1357_;
  (* src = "CanBsp.scala:270.117" *)
  wire _1358_;
  (* src = "CanBsp.scala:270.101" *)
  wire _1359_;
  (* src = "CanBsp.scala:270.82" *)
  wire _1360_;
  (* src = "Cat.scala:30.58" *)
  wire [8:0] _1361_;
  (* src = "CanBsp.scala:844.43" *)
  wire [9:0] _1362_;
  (* src = "CanBsp.scala:844.43" *)
  wire [8:0] _1363_;
  (* src = "CanBsp.scala:848.43" *)
  wire [9:0] _1364_;
  (* src = "CanBsp.scala:848.43" *)
  wire [8:0] _1365_;
  (* src = "CanBsp.scala:851.43" *)
  wire [9:0] _1366_;
  (* src = "CanBsp.scala:851.43" *)
  wire [8:0] _1367_;
  (* src = "CanBsp.scala:233.40" *)
  wire _1368_;
  (* src = "CanBsp.scala:233.56" *)
  wire _1369_;
  (* src = "CanBsp.scala:233.86" *)
  wire _1370_;
  (* src = "CanBsp.scala:795.30" *)
  wire [3:0] _1371_;
  (* src = "CanBsp.scala:795.30" *)
  wire [2:0] _1372_;
  (* src = "CanBsp.scala:407.27" *)
  wire [6:0] _1373_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _1374_;
  (* src = "CanBsp.scala:722.54" *)
  wire [63:0] _1375_;
  (* src = "CanBsp.scala:728.50" *)
  wire _1376_;
  (* src = "CanBsp.scala:728.78" *)
  wire [18:0] _1377_;
  (* src = "CanBsp.scala:728.78" *)
  wire _1378_;
  (* src = "CanBsp.scala:728.19" *)
  wire _1379_;
  (* src = "CanBsp.scala:732.30" *)
  wire [63:0] _1380_;
  (* src = "CanBsp.scala:732.30" *)
  wire _1381_;
  (* src = "CanBsp.scala:738.26" *)
  wire [18:0] _1382_;
  (* src = "CanBsp.scala:738.26" *)
  wire _1383_;
  (* src = "CanBsp.scala:722.54" *)
  wire _1384_;
  (* src = "CanBsp.scala:722.86" *)
  wire [63:0] _1385_;
  (* src = "CanBsp.scala:722.86" *)
  wire _1386_;
  (* src = "CanBsp.scala:722.19" *)
  wire _1387_;
  (* src = "CanBsp.scala:724.30" *)
  wire [14:0] _1388_;
  (* src = "CanBsp.scala:724.30" *)
  wire _1389_;
  (* src = "CanBsp.scala:728.50" *)
  wire [38:0] _1390_;
  (* src = "CanBsp.scala:863.36" *)
  wire [9:0] _1391_;
  (* src = "CanBsp.scala:863.36" *)
  wire [8:0] _1392_;
  (* src = "CanBsp.scala:869.38" *)
  wire [9:0] _1393_;
  (* src = "CanBsp.scala:869.38" *)
  wire [8:0] _1394_;
  (* src = "CanBsp.scala:111.36" *)
  wire _1395_;
  (* src = "CanBsp.scala:745.28" *)
  wire [6:0] _1396_;
  (* src = "CanBsp.scala:745.28" *)
  wire [5:0] _1397_;
  (* src = "CanBsp.scala:717.20" *)
  wire _1398_;
  (* src = "CanBsp.scala:717.18" *)
  wire _1399_;
  (* src = "CanBsp.scala:77.36" *)
  wire _1400_;
  wire [7:0] _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire [2:0] _1410_;
  wire _1411_;
  wire [2:0] _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire [2:0] _1416_;
  wire _1417_;
  wire [2:0] _1418_;
  wire _1419_;
  wire [2:0] _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire [2:0] _1426_;
  wire _1427_;
  wire [2:0] _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire [2:0] _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire [7:0] _1438_;
  wire _1439_;
  wire [14:0] _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire [2:0] _1480_;
  wire _1481_;
  wire [2:0] _1482_;
  wire _1483_;
  wire [28:0] _1484_;
  wire _1485_;
  wire [3:0] _1486_;
  wire _1487_;
  wire [5:0] _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire [4:0] _1494_;
  wire _1495_;
  wire [8:0] _1496_;
  wire _1497_;
  wire [8:0] _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire [7:0] _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire [2:0] _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire [3:0] _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire [5:0] _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire [4:0] _1562_;
  wire _1563_;
  (* src = "CanBsp.scala:232.75" *)
  wire ackErr;
  (* src = "CanBsp.scala:172.37" *)
  reg ackErrLatched;
  (* src = "CanBsp.scala:172.37|CanBsp.scala:172.37" *)
  wire \ackErrLatched$process$CanBsp_72 ;
  (* src = "CanBsp.scala:158.42" *)
  reg arbitrationBlocked;
  (* src = "CanBsp.scala:158.42|CanBsp.scala:158.42" *)
  wire \arbitrationBlocked$process$CanBsp_60 ;
  (* src = "CanBsp.scala:157.38" *)
  reg [4:0] arbitrationCnt;
  (* src = "CanBsp.scala:157.38|CanBsp.scala:157.38" *)
  wire [4:0] \arbitrationCnt$process$CanBsp_59 ;
  (* src = "CanBsp.scala:247.64" *)
  wire arbitrationField;
  (* src = "CanBsp.scala:156.41" *)
  reg arbitrationFieldD;
  (* src = "CanBsp.scala:156.41|CanBsp.scala:156.41" *)
  wire \arbitrationFieldD$process$CanBsp_58 ;
  (* src = "CanBsp.scala:154.39" *)
  reg arbitrationLost;
  (* src = "CanBsp.scala:154.39|CanBsp.scala:154.39" *)
  wire \arbitrationLost$process$CanBsp_56 ;
  (* src = "CanBsp.scala:99.46" *)
  reg [4:0] arbitrationLostCapture;
  (* src = "CanBsp.scala:99.46|CanBsp.scala:99.46" *)
  wire [4:0] \arbitrationLostCapture$process$CanBsp_11 ;
  (* src = "CanBsp.scala:155.40" *)
  reg arbitrationLostQ;
  (* src = "CanBsp.scala:155.40|CanBsp.scala:155.40|CanBsp.scala:155.40" *)
  wire \arbitrationLostQ$process$CanBsp_57 ;
  (* src = "Cat.scala:30.58" *)
  wire [18:0] basicChain;
  (* src = "Cat.scala:30.58" *)
  wire [63:0] basicChainData;
  (* src = "CanBsp.scala:106.30" *)
  reg [5:0] bitCnt;
  (* src = "CanBsp.scala:106.30|CanBsp.scala:106.30" *)
  wire [5:0] \bitCnt$process$CanBsp_15 ;
  (* src = "CanBsp.scala:188.39" *)
  wire bitDeStuff;
  (* src = "CanBsp.scala:215.58" *)
  wire bitDeStuffReset;
  (* src = "CanBsp.scala:214.38" *)
  wire bitDeStuffSet;
  (* src = "CanBsp.scala:189.43" *)
  wire bitDeStuffTx;
  (* src = "CanBsp.scala:269.207" *)
  wire bitErr;
  (* src = "CanBsp.scala:225.46" *)
  wire bitErrCompGoRxCrc;
  (* src = "CanBsp.scala:261.57" *)
  wire bitErrExc1;
  (* src = "CanBsp.scala:262.33" *)
  wire bitErrExc2;
  (* src = "CanBsp.scala:263.60" *)
  wire bitErrExc3;
  (* src = "CanBsp.scala:264.82" *)
  wire bitErrExc4;
  (* src = "CanBsp.scala:265.61" *)
  wire bitErrExc5;
  (* src = "CanBsp.scala:266.52" *)
  wire bitErrExc6;
  (* src = "CanBsp.scala:173.37" *)
  reg bitErrLatched;
  (* src = "CanBsp.scala:173.37|CanBsp.scala:173.37" *)
  wire \bitErrLatched$process$CanBsp_73 ;
  (* src = "CanBsp.scala:109.35" *)
  reg [2:0] bitStuffCnt;
  (* src = "CanBsp.scala:109.35|CanBsp.scala:109.35" *)
  wire [2:0] \bitStuffCnt$process$CanBsp_18 ;
  (* src = "CanBsp.scala:139.37" *)
  reg bitStuffCntEn;
  (* src = "CanBsp.scala:139.37|CanBsp.scala:139.37" *)
  wire \bitStuffCntEn$process$CanBsp_43 ;
  (* src = "CanBsp.scala:110.37" *)
  reg [2:0] bitStuffCntTx;
  (* src = "CanBsp.scala:110.37|CanBsp.scala:110.37" *)
  wire [2:0] \bitStuffCntTx$process$CanBsp_19 ;
  (* src = "CanBsp.scala:170.31" *)
  reg busFree;
  (* src = "CanBsp.scala:170.31|CanBsp.scala:170.31" *)
  wire \busFree$process$CanBsp_70 ;
  (* src = "CanBsp.scala:167.34" *)
  reg [3:0] busFreeCnt;
  (* src = "CanBsp.scala:167.34|CanBsp.scala:167.34" *)
  wire [3:0] \busFreeCnt$process$CanBsp_67 ;
  (* src = "CanBsp.scala:168.36" *)
  reg busFreeCntEn;
  (* src = "CanBsp.scala:168.36|CanBsp.scala:168.36" *)
  wire \busFreeCntEn$process$CanBsp_68 ;
  (* src = "CanBsp.scala:138.31" *)
  reg [2:0] byteCnt;
  (* src = "CanBsp.scala:138.31|CanBsp.scala:138.31" *)
  wire [2:0] \byteCnt$process$CanBsp_42 ;
  (* src = "CanBsp.scala:219.34|CanBsp.scala:524.17" *)
  wire [14:0] calculatedCrc;
  (* src = "CanBsp.scala:237.25|CanBsp.scala:543.8" *)
  wire canAcf_io_idOk;
  (* src = "CanBsp.scala:219.34|CanBsp.scala:524.17" *)
  wire [14:0] canCrcRx_io_crc;
  (* src = "CanBsp.scala:581.14" *)
  wire [7:0] canFifo_io_dataOut;
  (* src = "CanBsp.scala:586.23" *)
  wire [6:0] canFifo_io_infoCnt;
  (* src = "CanBsp.scala:587.16" *)
  wire canFifo_io_infoEmpty;
  (* src = "CanBsp.scala:585.14" *)
  wire canFifo_io_overrun;
  input clock;
  (* src = "CanBsp.scala:140.33" *)
  reg crcEnable;
  (* src = "CanBsp.scala:140.33|CanBsp.scala:140.33" *)
  wire \crcEnable$process$CanBsp_44 ;
  (* src = "CanBsp.scala:153.30" *)
  reg crcErr;
  (* src = "CanBsp.scala:153.30|CanBsp.scala:153.30" *)
  wire \crcErr$process$CanBsp_55 ;
  (* src = "CanBsp.scala:130.29" *)
  reg [14:0] crcIn;
  (* src = "CanBsp.scala:130.29|CanBsp.scala:130.29" *)
  wire [14:0] \crcIn$process$CanBsp_39 ;
  (* src = "CanBsp.scala:160.31" *)
  reg [3:0] dataCnt;
  (* src = "CanBsp.scala:160.31|CanBsp.scala:160.31" *)
  wire [3:0] \dataCnt$process$CanBsp_62 ;
  (* src = "CanBsp.scala:107.31" *)
  reg [3:0] dataLen;
  (* src = "CanBsp.scala:107.31|CanBsp.scala:107.31" *)
  wire [3:0] \dataLen$process$CanBsp_16 ;
  (* src = "CanBsp.scala:147.42" *)
  reg [2:0] delayedDominantCnt;
  (* src = "CanBsp.scala:147.42|CanBsp.scala:147.42" *)
  wire [2:0] \delayedDominantCnt$process$CanBsp_51 ;
  (* src = "CanBsp.scala:144.39" *)
  reg enableErrorCnt2;
  (* src = "CanBsp.scala:144.39|CanBsp.scala:144.39" *)
  wire \enableErrorCnt2$process$CanBsp_48 ;
  (* src = "CanBsp.scala:148.42" *)
  reg enableOverloadCnt2;
  (* src = "CanBsp.scala:148.42|CanBsp.scala:148.42" *)
  wire \enableOverloadCnt2$process$CanBsp_52 ;
  (* src = "CanBsp.scala:141.30" *)
  reg [2:0] eofCnt;
  (* src = "CanBsp.scala:141.30|CanBsp.scala:141.30" *)
  wire [2:0] \eofCnt$process$CanBsp_45 ;
  (* src = "CanBsp.scala:245.124" *)
  wire err;
  (* src = "CanBsp.scala:81.40" *)
  reg [7:0] errorCaptureCode;
  (* src = "CanBsp.scala:81.40|CanBsp.scala:81.40" *)
  wire [7:0] \errorCaptureCode$process$CanBsp_2 ;
  (* src = "CanBsp.scala:182.47" *)
  reg errorCaptureCodeBlocked;
  (* src = "CanBsp.scala:182.47|CanBsp.scala:182.47" *)
  wire \errorCaptureCodeBlocked$process$CanBsp_82 ;
  (* src = "CanBsp.scala:186.42" *)
  wire errorCaptureCodeDirection;
  (* src = "CanBsp.scala:925.16|CanBsp.scala:926.26" *)
  wire [1:0] errorCaptureCodeType;
  (* src = "CanBsp.scala:145.33" *)
  reg [2:0] errorCnt1;
  (* src = "CanBsp.scala:145.33|CanBsp.scala:145.33" *)
  wire [2:0] \errorCnt1$process$CanBsp_49 ;
  (* src = "CanBsp.scala:146.33" *)
  reg [2:0] errorCnt2;
  (* src = "CanBsp.scala:146.33|CanBsp.scala:146.33" *)
  wire [2:0] \errorCnt2$process$CanBsp_50 ;
  (* src = "CanBsp.scala:267.155" *)
  wire errorFlagOver;
  (* src = "CanBsp.scala:180.44" *)
  reg errorFlagOverLatched;
  (* src = "CanBsp.scala:180.44|CanBsp.scala:180.44" *)
  wire \errorFlagOverLatched$process$CanBsp_81 ;
  (* src = "CanBsp.scala:143.34" *)
  reg errorFrame;
  (* src = "CanBsp.scala:143.34|CanBsp.scala:143.34" *)
  wire \errorFrame$process$CanBsp_47 ;
  (* src = "CanBsp.scala:229.51" *)
  wire errorFrameEnded;
  (* src = "Cat.scala:30.58" *)
  wire [63:0] extendedChainDataExt;
  (* src = "Cat.scala:30.58" *)
  wire [63:0] extendedChainDataStd;
  (* src = "Cat.scala:30.58" *)
  wire [38:0] extendedChainExt;
  (* src = "Cat.scala:30.58" *)
  wire [18:0] extendedChainStd;
  (* src = "Cat.scala:30.58" *)
  wire [5:0] fifoSelector;
  (* src = "CanBsp.scala:166.33" *)
  reg finishMsg;
  (* src = "CanBsp.scala:166.33|CanBsp.scala:166.33" *)
  wire \finishMsg$process$CanBsp_66 ;
  (* src = "CanBsp.scala:183.39" *)
  reg firstCompareBit;
  (* src = "CanBsp.scala:183.39|CanBsp.scala:183.39" *)
  wire \firstCompareBit$process$CanBsp_83 ;
  (* src = "CanBsp.scala:222.39" *)
  wire formErr;
  (* src = "CanBsp.scala:175.38" *)
  reg formErrLatched;
  (* src = "CanBsp.scala:175.38|CanBsp.scala:175.38" *)
  wire \formErrLatched$process$CanBsp_75 ;
  (* src = "CanBsp.scala:211.40" *)
  wire goCrcEnable;
  (* src = "CanBsp.scala:217.149" *)
  wire goEarlyTx;
  (* src = "CanBsp.scala:126.40" *)
  reg goEarlyTxLatched;
  (* src = "CanBsp.scala:126.40|CanBsp.scala:126.40" *)
  wire \goEarlyTxLatched$process$CanBsp_35 ;
  (* src = "CanBsp.scala:206.55" *)
  wire goRxAck;
  (* src = "CanBsp.scala:207.42" *)
  wire goRxAckLim;
  (* src = "CanBsp.scala:227.45" *)
  wire goRxCrc;
  (* src = "CanBsp.scala:205.66" *)
  wire goRxCrcLim;
  (* src = "CanBsp.scala:226.117" *)
  wire goRxData;
  (* src = "CanBsp.scala:202.55" *)
  wire goRxDlc;
  (* src = "CanBsp.scala:208.39" *)
  wire goRxEof;
  (* src = "CanBsp.scala:195.56" *)
  wire goRxId1;
  (* src = "CanBsp.scala:198.63" *)
  wire goRxId2;
  (* src = "CanBsp.scala:197.55" *)
  wire goRxIde;
  (* src = "CanBsp.scala:194.73" *)
  wire goRxIdle;
  (* src = "CanBsp.scala:201.54" *)
  wire goRxR0;
  (* src = "CanBsp.scala:200.54" *)
  wire goRxR1;
  (* src = "CanBsp.scala:196.64" *)
  wire goRxRtr1;
  (* src = "CanBsp.scala:199.64" *)
  wire goRxRtr2;
  (* src = "CanBsp.scala:161.33" *)
  reg [2:0] headerCnt;
  (* src = "CanBsp.scala:161.33|CanBsp.scala:161.33" *)
  wire [2:0] \headerCnt$process$CanBsp_63 ;
  (* src = "CanBsp.scala:241.29" *)
  wire [2:0] headerLen;
  (* src = "CanBsp.scala:108.26" *)
  reg [28:0] id;
  (* src = "CanBsp.scala:108.26|CanBsp.scala:108.26" *)
  wire [28:0] \id$process$CanBsp_17 ;
  (* src = "CanBsp.scala:237.25|CanBsp.scala:543.8" *)
  wire idOk;
  (* src = "CanBsp.scala:128.27" *)
  reg ide;
  (* src = "CanBsp.scala:128.27|CanBsp.scala:128.27" *)
  wire \ide$process$CanBsp_37 ;
  input io_abortTx;
  input [7:0] io_acceptanceCode_0;
  input [7:0] io_acceptanceCode_1;
  input [7:0] io_acceptanceCode_2;
  input [7:0] io_acceptanceCode_3;
  input io_acceptanceFilterMode;
  input [7:0] io_acceptanceMask_0;
  input [7:0] io_acceptanceMask_1;
  input [7:0] io_acceptanceMask_2;
  input [7:0] io_acceptanceMask_3;
  input [7:0] io_addr;
  output [4:0] io_arbitrationLostCapture;
  output io_busOffOn;
  input [7:0] io_dataIn;
  output [7:0] io_dataOut;
  output [7:0] io_errorCaptureCode;
  output io_errorStatus;
  input [7:0] io_errorWarningLimit;
  input io_extendedMode;
  output io_goErrorFrame;
  output io_goOverloadFrame;
  output io_goRxInter;
  output io_goTx;
  input io_hardSync;
  output io_infoEmpty;
  input io_listenOnlyMode;
  output io_needToTx;
  output io_nodeBusOff;
  output io_nodeErrorActive;
  output io_nodeErrorPassive;
  output io_notFirstBitOfInter;
  output io_overloadFrame;
  output io_overrun;
  input io_readArbitrationLostCaptureReg;
  input io_readErrorCodeCaptureReg;
  output io_receiveStatus;
  input io_releaseBuffer;
  input io_resetMode;
  output [8:0] io_rxErrorCount;
  output io_rxIdle;
  output io_rxInter;
  output [6:0] io_rxMessageCounter;
  input io_samplePoint;
  input io_sampledBit;
  input io_sampledBitQ;
  input io_selfRxRequest;
  input io_selfTestMode;
  output io_sendAck;
  output io_setArbitrationLostIrq;
  output io_setBusErrorIrq;
  output io_setResetMode;
  input io_singleShotTransmission;
  output io_transmitStatus;
  output io_transmitter;
  output io_transmitting;
  output io_tx;
  input [7:0] io_txData_0;
  input [7:0] io_txData_1;
  input [7:0] io_txData_10;
  input [7:0] io_txData_11;
  input [7:0] io_txData_12;
  input [7:0] io_txData_2;
  input [7:0] io_txData_3;
  input [7:0] io_txData_4;
  input [7:0] io_txData_5;
  input [7:0] io_txData_6;
  input [7:0] io_txData_7;
  input [7:0] io_txData_8;
  input [7:0] io_txData_9;
  output [8:0] io_txErrorCount;
  output io_txNext;
  input io_txPoint;
  input io_txRequest;
  output io_txState;
  output io_txStateQ;
  output io_txSuccessful;
  input io_writeEnReceiveErrorCounter;
  input io_writeEnTransmitErrorCounter;
  (* src = "CanBsp.scala:192.39" *)
  wire lastBitOfInter;
  (* src = "CanBsp.scala:221.34" *)
  wire [3:0] limitedDataLen;
  (* src = "CanBsp.scala:243.40" *)
  wire [3:0] limitedDataLenSubOne;
  (* src = "CanBsp.scala:271.35" *)
  wire [5:0] limitedTxCntExt;
  (* src = "CanBsp.scala:272.35" *)
  wire [5:0] limitedTxCntStd;
  (* src = "CanBsp.scala:93.32" *)
  reg needToTx;
  (* src = "CanBsp.scala:93.32|CanBsp.scala:93.32" *)
  wire \needToTx$process$CanBsp_8 ;
  (* src = "CanBsp.scala:91.34" *)
  reg nodeBusOff;
  (* src = "CanBsp.scala:91.34|CanBsp.scala:91.34" *)
  wire \nodeBusOff$process$CanBsp_7 ;
  (* src = "CanBsp.scala:171.35" *)
  reg nodeBusOffQ;
  (* src = "CanBsp.scala:171.35|CanBsp.scala:171.35|CanBsp.scala:171.35" *)
  wire \nodeBusOffQ$process$CanBsp_71 ;
  (* src = "CanBsp.scala:101.40" *)
  reg nodeErrorPassive;
  (* src = "CanBsp.scala:101.40|CanBsp.scala:101.40" *)
  wire \nodeErrorPassive$process$CanBsp_12 ;
  (* src = "CanBsp.scala:151.36" *)
  reg [2:0] overloadCnt1;
  (* src = "CanBsp.scala:151.36|CanBsp.scala:151.36" *)
  wire [2:0] \overloadCnt1$process$CanBsp_53 ;
  (* src = "CanBsp.scala:152.36" *)
  reg [2:0] overloadCnt2;
  (* src = "CanBsp.scala:152.36|CanBsp.scala:152.36" *)
  wire [2:0] \overloadCnt2$process$CanBsp_54 ;
  (* src = "CanBsp.scala:268.73" *)
  wire overloadFlagOver;
  (* src = "CanBsp.scala:79.37" *)
  reg overloadFrame;
  (* src = "CanBsp.scala:79.37|CanBsp.scala:79.37" *)
  wire \overloadFrame$process$CanBsp_1 ;
  (* src = "CanBsp.scala:230.58" *)
  wire overloadFrameEnded;
  (* src = "CanBsp.scala:142.34" *)
  reg [2:0] passiveCnt;
  (* src = "CanBsp.scala:142.34|CanBsp.scala:142.34" *)
  wire [2:0] \passiveCnt$process$CanBsp_46 ;
  (* src = "Cat.scala:30.58" *)
  wire [14:0] rCalculatedCrc;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_0;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_1;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_10;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_11;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_12;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_2;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_3;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_4;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_5;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_6;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_7;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_8;
  (* src = "Bitwise.scala:103.39" *)
  wire [7:0] rTxData_9;
  (* src = "CanBsp.scala:209.41" *)
  wire remoteRq;
  input reset;
  (* src = "CanBsp.scala:105.34" *)
  reg resetModeQ;
  (* src = "CanBsp.scala:105.34|CanBsp.scala:105.34|CanBsp.scala:105.34" *)
  wire \resetModeQ$process$CanBsp_14 ;
  (* src = "CanBsp.scala:244.78" *)
  wire resetWrFifo;
  (* src = "CanBsp.scala:279.139" *)
  wire rstTxPointer;
  (* src = "CanBsp.scala:127.28" *)
  reg rtr1;
  (* src = "CanBsp.scala:127.28|CanBsp.scala:127.28" *)
  wire \rtr1$process$CanBsp_36 ;
  (* src = "CanBsp.scala:129.28" *)
  reg rtr2;
  (* src = "CanBsp.scala:129.28|CanBsp.scala:129.28" *)
  wire \rtr2$process$CanBsp_38 ;
  (* src = "CanBsp.scala:176.38" *)
  reg rule3Exc1_0;
  (* src = "CanBsp.scala:176.38|CanBsp.scala:176.38" *)
  wire \rule3Exc1_0$process$CanBsp_76 ;
  (* src = "CanBsp.scala:176.38" *)
  reg rule3Exc1_1;
  (* src = "CanBsp.scala:176.38|CanBsp.scala:176.38" *)
  wire \rule3Exc1_1$process$CanBsp_77 ;
  (* src = "CanBsp.scala:270.19" *)
  wire rule5;
  (* src = "CanBsp.scala:123.29" *)
  reg rxAck;
  (* src = "CanBsp.scala:123.29|CanBsp.scala:123.29" *)
  wire \rxAck$process$CanBsp_32 ;
  (* src = "CanBsp.scala:124.32" *)
  reg rxAckLim;
  (* src = "CanBsp.scala:124.32|CanBsp.scala:124.32" *)
  wire \rxAckLim$process$CanBsp_33 ;
  (* src = "CanBsp.scala:121.29" *)
  reg rxCrc;
  (* src = "CanBsp.scala:121.29|CanBsp.scala:121.29" *)
  wire \rxCrc$process$CanBsp_30 ;
  (* src = "CanBsp.scala:122.32" *)
  reg rxCrcLim;
  (* src = "CanBsp.scala:122.32|CanBsp.scala:122.32" *)
  wire \rxCrcLim$process$CanBsp_31 ;
  (* src = "CanBsp.scala:120.30" *)
  reg rxData;
  (* src = "CanBsp.scala:120.30|CanBsp.scala:120.30" *)
  wire \rxData$process$CanBsp_29 ;
  (* src = "CanBsp.scala:119.29" *)
  reg rxDlc;
  (* src = "CanBsp.scala:119.29|CanBsp.scala:119.29" *)
  wire \rxDlc$process$CanBsp_28 ;
  (* src = "CanBsp.scala:125.29" *)
  reg rxEof;
  (* src = "CanBsp.scala:125.29|CanBsp.scala:125.29" *)
  wire \rxEof$process$CanBsp_34 ;
  (* src = "CanBsp.scala:95.36" *)
  reg [8:0] rxErrorCount;
  (* src = "CanBsp.scala:95.36|CanBsp.scala:95.36" *)
  wire [8:0] \rxErrorCount$process$CanBsp_9 ;
  (* src = "CanBsp.scala:112.29" *)
  reg rxId1;
  (* src = "CanBsp.scala:112.29|CanBsp.scala:112.29" *)
  wire \rxId1$process$CanBsp_21 ;
  (* src = "CanBsp.scala:115.29" *)
  reg rxId2;
  (* src = "CanBsp.scala:115.29|CanBsp.scala:115.29" *)
  wire \rxId2$process$CanBsp_24 ;
  (* src = "CanBsp.scala:114.29" *)
  reg rxIde;
  (* src = "CanBsp.scala:114.29|CanBsp.scala:114.29" *)
  wire \rxIde$process$CanBsp_23 ;
  (* src = "CanBsp.scala:83.30" *)
  reg rxIdle;
  (* src = "CanBsp.scala:83.30|CanBsp.scala:83.30" *)
  wire \rxIdle$process$CanBsp_3 ;
  (* src = "CanBsp.scala:89.31" *)
  reg rxInter;
  (* src = "CanBsp.scala:89.31|CanBsp.scala:89.31" *)
  wire \rxInter$process$CanBsp_6 ;
  (* src = "CanBsp.scala:117.28" *)
  reg rxR0;
  (* src = "CanBsp.scala:117.28|CanBsp.scala:117.28" *)
  wire \rxR0$process$CanBsp_26 ;
  (* src = "CanBsp.scala:118.27" *)
  reg rxR1;
  (* src = "CanBsp.scala:118.27|CanBsp.scala:118.27" *)
  wire \rxR1$process$CanBsp_27 ;
  (* src = "CanBsp.scala:113.30" *)
  reg rxRtr1;
  (* src = "CanBsp.scala:113.30|CanBsp.scala:113.30" *)
  wire \rxRtr1$process$CanBsp_22 ;
  (* src = "CanBsp.scala:116.30" *)
  reg rxRtr2;
  (* src = "CanBsp.scala:116.30|CanBsp.scala:116.30" *)
  wire \rxRtr2$process$CanBsp_25 ;
  (* src = "CanBsp.scala:242.40" *)
  wire storingHeader;
  (* src = "CanBsp.scala:233.69" *)
  wire stuffErr;
  (* src = "CanBsp.scala:174.39" *)
  reg stuffErrLatched;
  (* src = "CanBsp.scala:174.39|CanBsp.scala:174.39" *)
  wire \stuffErrLatched$process$CanBsp_74 ;
  (* src = "CanBsp.scala:177.31" *)
  reg suspend;
  (* src = "CanBsp.scala:177.31|CanBsp.scala:177.31" *)
  wire \suspend$process$CanBsp_78 ;
  (* src = "CanBsp.scala:179.34" *)
  reg [2:0] suspendCnt;
  (* src = "CanBsp.scala:179.34|CanBsp.scala:179.34" *)
  wire [2:0] \suspendCnt$process$CanBsp_80 ;
  (* src = "CanBsp.scala:178.36" *)
  reg suspendCntEn;
  (* src = "CanBsp.scala:178.36|CanBsp.scala:178.36" *)
  wire \suspendCntEn$process$CanBsp_79 ;
  (* src = "CanBsp.scala:131.31" *)
  reg [7:0] tmpData;
  (* src = "CanBsp.scala:131.31|CanBsp.scala:131.31" *)
  wire [7:0] \tmpData$process$CanBsp_40 ;
  wire [7:0] tmpFifo_canAcf_io_data0_MPORT_data;
  wire [7:0] tmpFifo_canAcf_io_data1_MPORT_data;
  wire [7:0] tmpFifo_dataForFifo_MPORT_data;
  (* src = "CanBsp.scala:87.35" *)
  reg transmitter;
  (* src = "CanBsp.scala:87.35|CanBsp.scala:87.35" *)
  wire \transmitter$process$CanBsp_5 ;
  (* src = "CanBsp.scala:85.36" *)
  reg transmitting;
  (* src = "CanBsp.scala:85.36|CanBsp.scala:85.36" *)
  wire \transmitting$process$CanBsp_4 ;
  (* src = "CanBsp.scala:103.26" *)
  reg tx;
  (* src = "CanBsp.scala:103.26|CanBsp.scala:103.26" *)
  wire \tx$process$CanBsp_13 ;
  (* src = "CanBsp.scala:720.25" *)
  wire txBit;
  (* src = "CanBsp.scala:97.36" *)
  reg [8:0] txErrorCount;
  (* src = "CanBsp.scala:97.36|CanBsp.scala:97.36" *)
  wire [8:0] \txErrorCount$process$CanBsp_10 ;
  (* src = "CanBsp.scala:111.32" *)
  reg txPointQ;
  (* src = "CanBsp.scala:111.32|CanBsp.scala:111.32|CanBsp.scala:111.32" *)
  wire \txPointQ$process$CanBsp_20 ;
  (* src = "CanBsp.scala:164.33" *)
  reg [5:0] txPointer;
  (* src = "CanBsp.scala:164.33|CanBsp.scala:164.33" *)
  wire [5:0] \txPointer$process$CanBsp_65 ;
  (* src = "CanBsp.scala:159.27" *)
  reg txQ;
  (* src = "CanBsp.scala:159.27|CanBsp.scala:159.27" *)
  wire \txQ$process$CanBsp_61 ;
  (* src = "CanBsp.scala:75.31" *)
  reg txState;
  (* src = "CanBsp.scala:75.31|CanBsp.scala:75.31" *)
  wire \txState$process$CanBsp ;
  (* src = "CanBsp.scala:77.32" *)
  reg txStateQ;
  (* src = "CanBsp.scala:77.32|CanBsp.scala:77.32|CanBsp.scala:77.32" *)
  wire \txStateQ$process$CanBsp_0 ;
  (* src = "CanBsp.scala:169.41" *)
  reg waitingForBusFree;
  (* src = "CanBsp.scala:169.41|CanBsp.scala:169.41" *)
  wire \waitingForBusFree$process$CanBsp_69 ;
  (* src = "CanBsp.scala:162.30" *)
  reg wrFifo;
  (* src = "CanBsp.scala:162.30|CanBsp.scala:162.30" *)
  wire \wrFifo$process$CanBsp_64 ;
  (* src = "CanBsp.scala:137.42" *)
  reg writeDataToTmpFifo;
  (* src = "CanBsp.scala:137.42|CanBsp.scala:137.42" *)
  wire \writeDataToTmpFifo$process$CanBsp_41 ;
  reg [7:0] tmpFifo [7:0];
  initial begin
    tmpFifo[0] = 8'h00;
    tmpFifo[1] = 8'h00;
    tmpFifo[2] = 8'h00;
    tmpFifo[3] = 8'h00;
    tmpFifo[4] = 8'h00;
    tmpFifo[5] = 8'h00;
    tmpFifo[6] = 8'h00;
    tmpFifo[7] = 8'h00;
  end
  always @(posedge clock) begin
    if (_1401_[0])
      tmpFifo[byteCnt][0:0] <= tmpData[0];
    if (_1401_[1])
      tmpFifo[byteCnt][1:1] <= tmpData[1];
    if (_1401_[2])
      tmpFifo[byteCnt][2:2] <= tmpData[2];
    if (_1401_[3])
      tmpFifo[byteCnt][3:3] <= tmpData[3];
    if (_1401_[4])
      tmpFifo[byteCnt][4:4] <= tmpData[4];
    if (_1401_[5])
      tmpFifo[byteCnt][5:5] <= tmpData[5];
    if (_1401_[6])
      tmpFifo[byteCnt][6:6] <= tmpData[6];
    if (_1401_[7])
      tmpFifo[byteCnt][7:7] <= tmpData[7];
  end
  assign tmpFifo_dataForFifo_MPORT_data = tmpFifo[_0823_[2:0]];
  assign tmpFifo_canAcf_io_data1_MPORT_data = tmpFifo[3'h1];
  assign tmpFifo_canAcf_io_data0_MPORT_data = tmpFifo[3'h0];
  assign _1322_ = { 1'h0, limitedDataLenSubOne } + { 1'h0, _0097_ };
  assign _0807_ = { 1'h0, byteCnt } + 4'h1;
  assign _0756_ = { 1'h0, bitCnt } + 7'h01;
  assign _1064_ = { 1'h0, passiveCnt } + 4'h1;
  assign _1058_ = { 1'h0, overloadCnt1 } + 4'h1;
  assign _1060_ = { 1'h0, overloadCnt2 } + 4'h1;
  assign _1396_ = { 1'h0, txPointer } + 7'h01;
  assign _1371_ = { 1'h0, suspendCnt } + 4'h1;
  assign _0749_ = { 1'h0, arbitrationCnt } + 6'h01;
  assign _1364_ = { 1'h0, io_rxErrorCount } + 10'h001;
  assign _1366_ = { 1'h0, io_rxErrorCount } + 10'h008;
  assign _1393_ = { 1'h0, txErrorCount } + 10'h008;
  assign _0801_ = { 1'h0, busFreeCnt } + 5'h01;
  assign _0851_ = { 1'h0, eofCnt } + 4'h1;
  assign _0799_ = { 1'h0, bitStuffCnt } + 4'h1;
  assign _0797_ = { 1'h0, bitStuffCntTx } + 4'h1;
  assign _0982_ = { 1'h0, headerCnt } + 4'h1;
  assign _0813_ = { 1'h0, dataCnt } + 5'h01;
  assign _0908_ = { 1'h0, errorCnt1 } + 4'h1;
  assign _0910_ = { 1'h0, errorCnt2 } + 4'h1;
  assign _0849_ = { 1'h0, delayedDominantCnt } + 4'h1;
  assign _1401_ = $signed(writeDataToTmpFifo) & (* src = "CanBsp.scala:136.32" *) $signed(1'h1);
  assign _0803_ = io_samplePoint & io_sampledBit;
  assign _0805_ = _0803_ & _0804_;
  assign goRxRtr1 = _0976_ & _0978_;
  assign _1285_ = _1284_ & 8'hcc;
  assign _1289_ = _0106_ & 8'h55;
  assign _1292_ = _1291_ & 8'haa;
  assign _1294_ = _0107_ & 8'h0f;
  assign _1297_ = _1296_ & 8'hf0;
  assign _1301_ = _0108_ & 8'h33;
  assign _1304_ = _1303_ & 8'hcc;
  assign _1308_ = _0109_ & 8'h55;
  assign _1311_ = _1310_ & 8'haa;
  assign _1313_ = _0110_ & 8'h0f;
  assign goRxIde = _0975_ & rxRtr1;
  assign _1316_ = _1315_ & 8'hf0;
  assign _1098_ = _0111_ & 8'h33;
  assign _1101_ = _1100_ & 8'hcc;
  assign _1104_ = _0112_ & 8'h55;
  assign _1107_ = _1106_ & 8'haa;
  assign _1109_ = _0113_ & 8'h0f;
  assign _1113_ = _1112_ & 8'hf0;
  assign _1116_ = _0114_ & 8'h33;
  assign _1120_ = _1119_ & 8'hcc;
  assign _1123_ = _0116_ & 8'h55;
  assign _0968_ = _0975_ & rxIde;
  assign _1127_ = _1126_ & 8'haa;
  assign _1129_ = _0117_ & 8'h0f;
  assign _1133_ = _1132_ & 8'hf0;
  assign _1136_ = _0118_ & 8'h33;
  assign _1139_ = _1138_ & 8'hcc;
  assign _1142_ = _0119_ & 8'h55;
  assign _1146_ = _1145_ & 8'haa;
  assign _1148_ = _0120_ & 8'h0f;
  assign _1152_ = _1150_ & 8'hf0;
  assign _1155_ = _0121_ & 8'h33;
  assign goRxId2 = _0968_ & io_sampledBit;
  assign _1158_ = _1157_ & 8'hcc;
  assign _1161_ = _0122_ & 8'h55;
  assign _1165_ = _1163_ & 8'haa;
  assign _1167_ = _0123_ & 8'h0f;
  assign _1170_ = _1169_ & 8'hf0;
  assign _1173_ = _0124_ & 8'h33;
  assign _1177_ = _1175_ & 8'hcc;
  assign _1180_ = _0125_ & 8'h55;
  assign _1184_ = _1182_ & 8'haa;
  assign _1186_ = _0127_ & 8'h0f;
  assign _0979_ = _0975_ & rxId2;
  assign _1189_ = _1188_ & 8'hf0;
  assign _1193_ = _0128_ & 8'h33;
  assign _1196_ = _1195_ & 8'hcc;
  assign _1200_ = _0129_ & 8'h55;
  assign _1203_ = _1202_ & 8'haa;
  assign _1205_ = _0130_ & 8'h0f;
  assign _1208_ = _1207_ & 8'hf0;
  assign _1212_ = _0131_ & 8'h33;
  assign _1215_ = _1214_ & 8'hcc;
  assign _1218_ = _0132_ & 8'h55;
  assign goRxRtr2 = _0979_ & _0981_;
  assign _1221_ = _1220_ & 8'haa;
  assign _1223_ = _0133_ & 8'h0f;
  assign _1226_ = _1225_ & 8'hf0;
  assign _1230_ = _0134_ & 8'h33;
  assign _1233_ = _1232_ & 8'hcc;
  assign _1237_ = _0135_ & 8'h55;
  assign _1240_ = _1239_ & 8'haa;
  assign _1243_ = _0136_ & 8'h0f;
  assign _1246_ = _1245_ & 8'hf0;
  assign _1250_ = _0138_ & 8'h33;
  assign goRxR1 = _0975_ & rxRtr2;
  assign _1253_ = _1252_ & 8'hcc;
  assign _1257_ = _0139_ & 8'h55;
  assign _1260_ = _1259_ & 8'haa;
  assign _1262_ = _0140_ & 8'h0f;
  assign _1265_ = _1264_ & 8'hf0;
  assign _1269_ = _0141_ & 8'h33;
  assign _1272_ = _1271_ & 8'hcc;
  assign _1276_ = _0142_ & 8'h55;
  assign _1279_ = _1278_ & 8'haa;
  assign _1020_ = _0941_ & rxAck;
  assign _0972_ = rxIde & _0965_;
  assign _1022_ = _1020_ & _1021_;
  assign _0913_ = _0912_ & io_samplePoint;
  assign _0914_ = _0913_ & _0767_;
  assign _0915_ = io_nodeErrorPassive & io_samplePoint;
  assign _0917_ = _0915_ & _0916_;
  assign errorFlagOver = _0918_ & _0769_;
  assign _1062_ = io_samplePoint & _0771_;
  assign overloadFlagOver = _1062_ & _0773_;
  assign _1356_ = _0912_ & errorFrame;
  assign _1357_ = _1356_ & _0766_;
  assign goRxR0 = _0975_ & _0973_;
  assign _1359_ = io_overloadFrame & _1358_;
  assign rule5 = bitErr & _1360_;
  assign _1325_ = _1324_ & io_txPoint;
  assign _1336_ = _1325_ & _1331_;
  assign _1342_ = _1336_ & io_extendedMode;
  assign _1353_ = _1342_ & _1352_;
  assign _1355_ = _1353_ & _1354_;
  assign _1327_ = _1342_ & _1326_;
  assign _1329_ = _1327_ & _1328_;
  assign _1333_ = _1336_ & _1332_;
  assign goRxDlc = _0975_ & rxR0;
  assign _1334_ = _1333_ & _1328_;
  assign _1337_ = _1325_ & rxData;
  assign _1338_ = _1337_ & io_extendedMode;
  assign _1340_ = _1338_ & _1339_;
  assign _1343_ = _1337_ & _1332_;
  assign _1345_ = _1343_ & _1344_;
  assign _1347_ = io_txPoint & rxCrcLim;
  assign _0999_ = rxEof & _0927_;
  assign _1000_ = _0999_ & _1005_;
  assign _1003_ = _0966_ & _1002_;
  assign _0806_ = _0805_ & waitingForBusFree;
  assign _0948_ = _0975_ & rxCrc;
  assign _0993_ = _0966_ & io_rxInter;
  assign _0995_ = _0993_ & _0994_;
  assign _0998_ = _0966_ & _0997_;
  assign _0992_ = crcErr & goRxEof;
  assign _1033_ = transmitter & io_goRxInter;
  assign _1034_ = _1033_ & _0759_;
  assign _1036_ = _1034_ & _1035_;
  assign _1038_ = _1036_ & _1037_;
  assign _0629_ = io_samplePoint & _0621_;
  assign _0646_ = _0629_ & _0974_;
  assign goRxCrcLim = _0948_ & _0949_;
  assign _0651_ = io_samplePoint & rxRtr1;
  assign _0669_ = _0651_ & _0974_;
  assign _0677_ = io_samplePoint & rxRtr2;
  assign _0693_ = _0677_ & _0974_;
  assign _0695_ = io_samplePoint & rxIde;
  assign _0696_ = _0695_ & _0974_;
  assign _0697_ = io_samplePoint & rxDlc;
  assign _0698_ = _0697_ & _0974_;
  assign _0699_ = io_samplePoint & rxData;
  assign _0700_ = _0699_ & _0974_;
  assign goRxAck = _0975_ & rxCrcLim;
  assign _0704_ = _0700_ & _0703_;
  assign _0705_ = io_samplePoint & goRxCrcLim;
  assign _0706_ = io_samplePoint & rxCrc;
  assign _0707_ = _0706_ & _0974_;
  assign _0719_ = io_samplePoint & _0974_;
  assign _0721_ = txPointQ & bitStuffCntEn;
  assign _0727_ = rule3Exc1_0 & _0766_;
  assign _0728_ = _0727_ & io_samplePoint;
  assign _0730_ = _0728_ & _0965_;
  assign _0732_ = io_transmitter & io_nodeErrorPassive;
  assign goRxAckLim = io_samplePoint & rxAck;
  assign _0733_ = _0732_ & ackErr;
  assign _0809_ = crcEnable & io_samplePoint;
  assign _0734_ = io_goRxInter & idOk;
  assign _0736_ = _0734_ & _1035_;
  assign _0738_ = _0736_ & _0737_;
  assign _0739_ = wrFifo & storingHeader;
  assign _0821_ = fifoSelector & 6'h37;
  assign _0744_ = errorFrame & io_txPoint;
  assign _0547_ = _0744_ & _0766_;
  assign _0548_ = errorFlagOver & io_sampledBit;
  assign goRxEof = io_samplePoint & rxAckLim;
  assign _0549_ = errorFrame & _0548_;
  assign _0551_ = enableErrorCnt2 & io_txPoint;
  assign _0556_ = _0966_ & _0555_;
  assign _0560_ = io_samplePoint & _0559_;
  assign _0561_ = errorFrame & _0769_;
  assign _0562_ = _0561_ & _1370_;
  assign _0565_ = io_overloadFrame & io_txPoint;
  assign _0566_ = _0565_ & _1358_;
  assign _0567_ = overloadFlagOver & io_sampledBit;
  assign _0568_ = io_overloadFrame & _0567_;
  assign _1320_ = _1319_ & rtr1;
  assign _0570_ = enableOverloadCnt2 & io_txPoint;
  assign _1029_ = _1324_ & txBit;
  assign _1031_ = bitDeStuffTx & _1030_;
  assign _1399_ = io_tx & _1398_;
  assign _0578_ = io_txPoint & _0577_;
  assign _0579_ = _0578_ & _1324_;
  assign _0583_ = io_abortTx & errorCaptureCodeDirection;
  assign _0585_ = _0941_ & io_txStateQ;
  assign _0586_ = _0585_ & io_singleShotTransmission;
  assign _0588_ = io_txRequest & io_samplePoint;
  assign _1321_ = ide & rtr2;
  assign _1008_ = io_samplePoint & _0944_;
  assign _1010_ = _0942_ & _1009_;
  assign _0595_ = suspend & goRxId1;
  assign _0601_ = goRxId1 & _0941_;
  assign _0603_ = arbitrationLost & io_txState;
  assign _0606_ = io_notFirstBitOfInter & io_transmitter;
  assign _0607_ = _0606_ & io_nodeErrorPassive;
  assign _0609_ = suspend & io_samplePoint;
  assign _0610_ = _0609_ & lastBitOfInter;
  assign _0611_ = suspendCntEn & io_samplePoint;
  assign bitDeStuffSet = goRxId1 & _0759_;
  assign _0617_ = io_transmitter & io_samplePoint;
  assign _0618_ = _0617_ & io_tx;
  assign _0619_ = _0618_ & arbitrationField;
  assign _0620_ = _0619_ & _0965_;
  assign _1024_ = arbitrationLost & _1023_;
  assign _0622_ = io_writeEnReceiveErrorCounter & _0970_;
  assign _0624_ = _0938_ & _0623_;
  assign _0625_ = goRxAckLim & _0759_;
  assign _0627_ = _0625_ & _0626_;
  assign _0630_ = _0627_ & _0628_;
  assign _0939_ = _0938_ & io_needToTx;
  assign _0634_ = io_goErrorFrame & _0633_;
  assign _0636_ = errorFlagOver & _0635_;
  assign _0637_ = _0636_ & io_samplePoint;
  assign _0638_ = _0637_ & _0965_;
  assign _0639_ = _0638_ & _0767_;
  assign _0640_ = io_goErrorFrame & rule5;
  assign _0643_ = _0966_ & _0642_;
  assign _0648_ = _0645_ & _0647_;
  assign _0649_ = io_transmitter & _1039_;
  assign _0653_ = io_goErrorFrame & _0652_;
  assign _0942_ = _0939_ & _0941_;
  assign _0654_ = io_transmitter & stuffErr;
  assign _0655_ = _0654_ & arbitrationField;
  assign _0656_ = _0655_ & io_samplePoint;
  assign _0657_ = _0656_ & io_tx;
  assign _0658_ = _0657_ & _0965_;
  assign _0660_ = _0653_ & _0659_;
  assign _0662_ = errorFrame & rule3Exc1_1;
  assign _0666_ = _0664_ & _0665_;
  assign _0671_ = _0788_ & resetModeQ;
  assign _0673_ = _0670_ & _0672_;
  assign lastBitOfInter = rxInter & _1041_;
  assign _0946_ = _0942_ & _0945_;
  assign _0674_ = _0673_ & _0970_;
  assign _0678_ = _0675_ & _0676_;
  assign _0679_ = _0678_ & _0788_;
  assign _0681_ = io_writeEnTransmitErrorCounter & _0680_;
  assign _0685_ = io_writeEnTransmitErrorCounter & _0684_;
  assign _0687_ = io_sampledBit & busFreeCntEn;
  assign _0689_ = _0687_ & _0688_;
  assign _0690_ = nodeBusOffQ & _0788_;
  assign _0694_ = _0805_ & _0970_;
  assign _0904_ = rxId2 & _0903_;
  assign _0947_ = _0946_ & io_samplePoint;
  assign _0873_ = rxId1 & _0871_;
  assign _0893_ = rxId2 & _0891_;
  assign _0900_ = errorFrame & io_nodeErrorActive;
  assign _1028_ = io_extendedMode & waitingForBusFree;
  assign _1015_ = _1014_ & errorCaptureCodeDirection;
  assign _1018_ = _1017_ & _1014_;
  assign _1019_ = _1018_ & errorCaptureCodeDirection;
  assign io_notFirstBitOfInter = io_rxInter & _1013_;
  assign io_setResetMode = nodeBusOff & _1027_;
  assign io_txSuccessful = _1038_ & _1039_;
  assign _0940_ = _0947_ & _0965_;
  assign io_setBusErrorIrq = io_goErrorFrame & _1026_;
  assign io_setArbitrationLostIrq = _1024_ & _1025_;
  assign io_goTx = _1010_ & _1011_;
  assign io_sendAck = _1022_ & _0938_;
  assign _0465_ = _0809_ & _0974_;
  assign _0466_ = _0948_ & _0949_;
  assign goEarlyTx = _0940_ & _0967_;
  assign _1088_ = _0094_ & 8'h0f;
  assign _1096_ = _1095_ & 8'hf0;
  assign _1068_ = _0095_ & 8'h33;
  assign _1071_ = _1070_ & 8'hcc;
  assign _1074_ = _0096_ & 8'h55;
  assign _1077_ = _1076_ & 8'haa;
  assign _0969_ = _0803_ & lastBitOfInter;
  assign _0925_ = _0974_ & rxCrcLim;
  assign _0933_ = _0925_ & _0965_;
  assign _0934_ = rxAckLim & _0965_;
  assign _0937_ = _0936_ & rxEof;
  assign _0926_ = _0937_ & _0965_;
  assign _0928_ = _0926_ & _0927_;
  assign _0930_ = rxEof & _0965_;
  assign _0931_ = _0930_ & io_transmitter;
  assign formErr = io_samplePoint & _0932_;
  assign _0958_ = _0975_ & rxDlc;
  assign _0971_ = busFree & _0970_;
  assign _0960_ = _0958_ & _0959_;
  assign _0964_ = _0960_ & _0963_;
  assign goRxData = _0964_ & _0957_;
  assign _0954_ = rxDlc & _0959_;
  assign _0956_ = _0965_ & _0955_;
  assign _0951_ = _0954_ & _0950_;
  assign _0952_ = rxData & bitErrCompGoRxCrc;
  assign goRxCrc = _0975_ & _0953_;
  assign errorFrameEnded = _0919_ & io_txPoint;
  assign overloadFrameEnded = _1063_ & io_txPoint;
  assign _0966_ = io_samplePoint & _0965_;
  assign _0745_ = rxAck & io_samplePoint;
  assign _0746_ = _0745_ & io_sampledBit;
  assign _0747_ = _0746_ & io_txState;
  assign ackErr = _0747_ & _0748_;
  assign _1368_ = io_samplePoint & bitStuffCntEn;
  assign _1369_ = _1368_ & bitDeStuff;
  assign stuffErr = _1369_ & _1370_;
  assign _1004_ = io_samplePoint & rxEof;
  assign _1006_ = _1004_ & _1005_;
  assign _0790_ = _0789_ & io_samplePoint;
  assign goRxId1 = _0966_ & _0967_;
  assign _0792_ = _0790_ & _0791_;
  assign _0764_ = io_txState & arbitrationField;
  assign bitErrExc1 = _0764_ & io_tx;
  assign _0794_ = _0792_ & _0793_;
  assign bitErrExc2 = rxAck & io_tx;
  assign _0796_ = _0794_ & _0795_;
  assign _0765_ = errorFrame & io_nodeErrorPassive;
  assign bitErrExc3 = _0765_ & _0766_;
  assign _0781_ = _0796_ & _0780_;
  assign _0768_ = errorFrame & _0767_;
  assign _0975_ = _0974_ & io_samplePoint;
  assign _0770_ = _0768_ & _0769_;
  assign _0772_ = io_overloadFrame & _0771_;
  assign _0774_ = _0772_ & _0773_;
  assign _0783_ = _0781_ & _0782_;
  assign _0775_ = errorFrame & _0919_;
  assign _0776_ = io_overloadFrame & _1063_;
  assign _0785_ = _0783_ & _0784_;
  assign _0777_ = _1005_ & rxEof;
  assign bitErrExc6 = _0777_ & _0927_;
  assign _0787_ = _0785_ & _0786_;
  assign _0976_ = _0975_ & rxId1;
  assign bitErr = _0787_ & _0788_;
  assign _1228_ = _0099_ & 8'h0f;
  assign _1299_ = _1287_ & 8'hf0;
  assign _1117_ = _0100_ & 8'h33;
  assign _1144_ = _1131_ & 8'hcc;
  assign _1183_ = _0101_ & 8'h55;
  assign _1210_ = _1197_ & 8'haa;
  assign _1241_ = _0102_ & 8'h0f;
  assign _1267_ = _1255_ & 8'hf0;
  assign _1282_ = _0105_ & 8'h33;
  assign _0804_ = busFreeCnt == 4'ha;
  assign bitDeStuff = bitStuffCnt == 3'h5;
  assign bitDeStuffTx = bitStuffCntTx == 3'h5;
  assign _1370_ = io_sampledBit == io_sampledBitQ;
  assign _1005_ = eofCnt == 3'h6;
  assign _1323_ = _0098_ == _1322_;
  assign _0771_ = overloadCnt1 == 3'h7;
  assign _0916_ = passiveCnt == 3'h6;
  assign _1354_ = txPointer == 6'h26;
  assign _1328_ = txPointer == 6'h12;
  assign _1339_ = txPointer == limitedTxCntExt;
  assign _1344_ = txPointer == limitedTxCntStd;
  assign _0722_ = io_tx == txQ;
  assign _1041_ = _1040_ == 2'h2;
  assign _0822_ = 6'h21 == _0821_;
  assign _0824_ = 6'h20 == _0821_;
  assign _0825_ = 6'h32 == fifoSelector;
  assign _0826_ = 6'h31 == fifoSelector;
  assign _0827_ = 6'h30 == fifoSelector;
  assign _0828_ = 6'h3c == fifoSelector;
  assign _0829_ = 6'h3b == fifoSelector;
  assign _0830_ = 6'h3a == fifoSelector;
  assign _0831_ = 6'h39 == fifoSelector;
  assign _0832_ = 6'h38 == fifoSelector;
  assign _0978_ = _0977_ == 4'ha;
  assign _0642_ = delayedDominantCnt == 3'h7;
  assign _0675_ = ! io_rxErrorCount;
  assign _0676_ = ! io_txErrorCount;
  assign _0684_ = io_dataIn == 8'hff;
  assign _0981_ = _0980_ == 5'h11;
  assign _0949_ = _0977_ == 4'he;
  assign _0944_ = suspendCnt == 3'h7;
  assign bitErrCompGoRxCrc = bitCnt == _0763_;
  assign _0959_ = _1040_ == 2'h3;
  assign _1063_ = overloadCnt2 == 3'h7;
  assign _0667_ = rxErrorCount >= 9'h080;
  assign _0668_ = txErrorCount >= 9'h080;
  assign _0683_ = io_txErrorCount >= 9'h100;
  assign _0986_ = io_rxErrorCount >= _0143_;
  assign _0987_ = io_txErrorCount >= _0143_;
  assign _0989_ = io_rxErrorCount >= 9'h060;
  assign _0990_ = io_txErrorCount >= 9'h060;
  assign _0628_ = io_rxErrorCount > 9'h000;
  assign _0631_ = io_rxErrorCount > 9'h07f;
  assign _0645_ = txErrorCount > 9'h000;
  assign _0903_ = bitCnt > 6'h04;
  assign _0871_ = bitCnt > 6'h07;
  assign _1045_ = dataLen < 4'h8;
  assign _0936_ = eofCnt < 3'h6;
  assign _1056_ = dataLen < 4'h1;
  assign _0632_ = io_rxErrorCount < 9'h080;
  assign _0664_ = rxErrorCount < 9'h080;
  assign _0665_ = txErrorCount < 9'h080;
  assign _0680_ = io_dataIn < 8'hff;
  assign _0688_ = busFreeCnt < 4'ha;
  assign _0891_ = bitCnt < 6'h0d;
  assign _1057_ = dataLen < 4'h2;
  assign storingHeader = headerCnt < headerLen;
  assign _0766_ = errorCnt1 < 3'h7;
  assign _1358_ = overloadCnt1 < 3'h7;
  assign _0994_ = _1040_ < 2'h2;
  assign _0559_ = passiveCnt < 3'h6;
  assign _0573_ = errorCnt1 < 3'h6;
  assign _0575_ = overloadCnt1 < 3'h6;
  assign _1400_ = io_resetMode ? (* src = "CanBsp.scala:77.36" *) 1'h0 : txState;
  assign _1395_ = io_resetMode ? (* src = "CanBsp.scala:111.36" *) 1'h0 : io_txPoint;
  assign limitedDataLen = _1045_ ? (* src = "CanBsp.scala:221.34" *) dataLen : 4'h8;
  assign _0168_ = _0613_ ? (* src = "CanBsp.scala:302.35|CanBsp.scala:303.12" *) 1'h0 : _0162_;
  assign _0017_ = _0574_ ? (* src = "CanBsp.scala:692.55" *) _0014_ : _0016_;
  assign _0018_ = _0206_ ? (* src = "CanBsp.scala:681.41" *) _0013_ : _0017_;
  assign _0020_ = io_txPoint ? (* src = "CanBsp.scala:710.26|CanBsp.scala:711.8|CanBsp.scala:103.26" *) io_txNext : tx;
  assign _0022_ = io_txPoint ? (* src = "CanBsp.scala:716.26|CanBsp.scala:717.9|CanBsp.scala:159.27" *) _1399_ : txQ;
  assign _0023_ = io_resetMode ? (* src = "CanBsp.scala:714.22|CanBsp.scala:715.9" *) 1'h0 : _0022_;
  assign _0031_ = _0580_ ? (* src = "CanBsp.scala:744.81|CanBsp.scala:745.15|CanBsp.scala:164.33" *) _1397_ : txPointer;
  assign _0032_ = rstTxPointer ? (* src = "CanBsp.scala:742.22|CanBsp.scala:743.15" *) 6'h00 : _0031_;
  assign _0034_ = _0587_ ? (* src = "CanBsp.scala:748.130|CanBsp.scala:749.14" *) 1'h0 : _0033_;
  assign _0036_ = _0589_ ? (* src = "CanBsp.scala:756.35|CanBsp.scala:757.22" *) 1'h0 : _0035_;
  assign _0038_ = _0593_ ? (* src = "CanBsp.scala:762.68|CanBsp.scala:763.13" *) 1'h0 : _0037_;
  assign _0190_ = _0701_ ? (* src = "CanBsp.scala:308.45|CanBsp.scala:309.11" *) 1'h0 : _0179_;
  assign _0040_ = _0596_ ? (* src = "CanBsp.scala:770.59|CanBsp.scala:771.17|CanBsp.scala:87.35" *) 1'h0 : transmitter;
  assign _0042_ = _0604_ ? (* src = "CanBsp.scala:776.98|CanBsp.scala:777.18|CanBsp.scala:85.36" *) 1'h0 : transmitting;
  assign _0045_ = _0605_ ? (* src = "CanBsp.scala:780.63|CanBsp.scala:781.13" *) 1'h0 : _0044_;
  assign _0047_ = _0605_ ? (* src = "CanBsp.scala:786.64|CanBsp.scala:787.18" *) 1'h0 : _0046_;
  assign _0048_ = _0611_ ? (* src = "CanBsp.scala:794.45|CanBsp.scala:795.16|CanBsp.scala:179.34" *) _1372_ : suspendCnt;
  assign _0049_ = _0605_ ? (* src = "CanBsp.scala:792.64|CanBsp.scala:793.16" *) 3'h0 : _0048_;
  assign _0052_ = _0615_ ? (* src = "CanBsp.scala:798.56|CanBsp.scala:799.15" *) 1'h0 : _0051_;
  assign _0054_ = _0616_ ? (* src = "CanBsp.scala:804.36|CanBsp.scala:805.21" *) 1'h0 : _0053_;
  assign _0055_ = io_samplePoint ? (* src = "CanBsp.scala:810.24|CanBsp.scala:811.23|CanBsp.scala:156.41" *) arbitrationField : arbitrationFieldD;
  assign _0056_ = arbitrationFieldD ? (* src = "CanBsp.scala:817.29|CanBsp.scala:818.22|CanBsp.scala:820.22" *) _0750_ : 5'h00;
  assign _0212_ = _0708_ ? (* src = "CanBsp.scala:314.37|CanBsp.scala:315.11" *) 1'h0 : _0201_;
  assign _0057_ = _0719_ ? (* src = "CanBsp.scala:816.38|CanBsp.scala:157.38" *) _0056_ : arbitrationCnt;
  assign _0058_ = io_setArbitrationLostIrq ? (* src = "CanBsp.scala:824.34|CanBsp.scala:825.28|CanBsp.scala:99.46" *) arbitrationCnt : arbitrationLostCapture;
  assign _0060_ = io_readArbitrationLostCaptureReg ? (* src = "CanBsp.scala:828.42|CanBsp.scala:829.24" *) 1'h0 : _0059_;
  assign _0062_ = _0631_ ? (* src = "CanBsp.scala:841.39|CanBsp.scala:842.24|CanBsp.scala:844.24" *) 9'h07f : _1363_;
  assign _0063_ = _0644_ ? (* src = "CanBsp.scala:850.116|CanBsp.scala:851.24|CanBsp.scala:95.36" *) _1367_ : rxErrorCount;
  assign _0064_ = _0634_ ? (* src = "CanBsp.scala:847.40|CanBsp.scala:848.24" *) _1365_ : _0063_;
  assign _0065_ = _0632_ ? (* src = "CanBsp.scala:846.43|CanBsp.scala:95.36" *) _0064_ : rxErrorCount;
  assign _0066_ = _0630_ ? (* src = "CanBsp.scala:840.83" *) _0062_ : _0065_;
  assign _0067_ = _0624_ ? (* src = "CanBsp.scala:839.68|CanBsp.scala:95.36" *) _0066_ : rxErrorCount;
  assign _0068_ = io_setResetMode ? (* src = "CanBsp.scala:836.30|CanBsp.scala:837.18" *) 9'h000 : _0067_;
  assign _0012_ = _0718_ ? (* src = "CanBsp.scala:320.34|CanBsp.scala:321.12" *) 1'h0 : _0002_;
  assign _0069_ = _0622_ ? (* src = "CanBsp.scala:834.58|CanBsp.scala:835.18" *) _1361_ : _0068_;
  assign _0070_ = _0663_ ? (* src = "CanBsp.scala:868.38|CanBsp.scala:869.22|CanBsp.scala:97.36" *) _1394_ : txErrorCount;
  assign _0071_ = _0649_ ? (* src = "CanBsp.scala:864.53|CanBsp.scala:97.36" *) _0070_ : txErrorCount;
  assign _0073_ = _0648_ ? (* src = "CanBsp.scala:862.68|CanBsp.scala:863.20" *) _1392_ : _0071_;
  assign _0074_ = io_setResetMode ? (* src = "CanBsp.scala:860.27|CanBsp.scala:861.20" *) 9'h080 : _0073_;
  assign _0075_ = io_writeEnTransmitErrorCounter ? (* src = "CanBsp.scala:857.40|CanBsp.scala:858.18" *) _1361_ : _0074_;
  assign _0077_ = _0666_ ? (* src = "CanBsp.scala:874.57|CanBsp.scala:875.22" *) 1'h0 : _0076_;
  assign _0079_ = _0682_ ? (* src = "CanBsp.scala:882.138|CanBsp.scala:883.16" *) 1'h0 : _0078_;
  assign _0080_ = _0689_ ? (* src = "CanBsp.scala:889.60|CanBsp.scala:890.18|CanBsp.scala:892.18" *) _0802_ : 4'h0;
  assign _0081_ = io_samplePoint ? (* src = "CanBsp.scala:888.24|CanBsp.scala:167.34" *) _0080_ : busFreeCnt;
  assign _0029_ = _0723_ ? (* src = "CanBsp.scala:326.34|CanBsp.scala:327.10" *) 1'h0 : _0019_;
  assign _0082_ = _0694_ ? (* src = "CanBsp.scala:898.87|CanBsp.scala:899.18|CanBsp.scala:168.36" *) 1'h0 : busFreeCntEn;
  assign _0086_ = _0971_ ? (* src = "CanBsp.scala:908.34|CanBsp.scala:909.23" *) 1'h0 : _0085_;
  assign _0089_ = stuffErr ? (* src = "CanBsp.scala:929.24|CanBsp.scala:930.26|CanBsp.scala:932.26" *) 2'h2 : 2'h3;
  assign _0090_ = formErr ? (* src = "CanBsp.scala:927.23|CanBsp.scala:928.26" *) 2'h1 : _0089_;
  assign errorCaptureCodeType = bitErr ? (* src = "CanBsp.scala:925.16|CanBsp.scala:926.26" *) 2'h0 : _0090_;
  assign _0087_ = io_setBusErrorIrq ? (* src = "CanBsp.scala:916.33|CanBsp.scala:917.22|CanBsp.scala:81.40" *) _0907_ : errorCaptureCode;
  assign _0088_ = io_readErrorCodeCaptureReg ? (* src = "CanBsp.scala:914.36|CanBsp.scala:915.22" *) 8'h00 : _0087_;
  assign _0093_ = io_readErrorCodeCaptureReg ? (* src = "CanBsp.scala:940.36|CanBsp.scala:941.29" *) 1'h0 : _0091_;
  assign _0144_ = reset ? (* src = "CanBsp.scala:160.31|CanBsp.scala:160.31" *) 5'h00 : _0205_;
  assign _0145_ = reset ? (* src = "CanBsp.scala:161.33|CanBsp.scala:161.33" *) 4'h0 : _0203_;
  assign _0050_ = _0729_ ? (* src = "CanBsp.scala:332.35|CanBsp.scala:333.10" *) 1'h0 : _0039_;
  assign io_errorStatus = io_extendedMode ? (* src = "CanBsp.scala:946.24" *) _0988_ : _0991_;
  assign io_receiveStatus = io_extendedMode ? (* src = "CanBsp.scala:936.27" *) _1016_ : _1019_;
  assign _0224_ = _0822_ ? (* src = "Lookup.scala:33.37" *) _0820_ : _0842_;
  assign _0072_ = _0546_ ? (* src = "CanBsp.scala:338.46|CanBsp.scala:339.11" *) 1'h0 : _0061_;
  assign _0092_ = _0550_ ? (* src = "CanBsp.scala:344.35|CanBsp.scala:345.12" *) 1'h0 : _0083_;
  assign _0115_ = _0557_ ? (* src = "CanBsp.scala:350.38|CanBsp.scala:351.11" *) 1'h0 : _0104_;
  assign _0137_ = _0758_ ? (* src = "CanBsp.scala:356.35|CanBsp.scala:357.14" *) 1'h0 : _0126_;
  assign _0983_ = ide ? (* src = "CanBsp.scala:241.50" *) 3'h5 : 3'h3;
  assign _0147_ = _0569_ ? (* src = "CanBsp.scala:362.38|CanBsp.scala:363.11" *) 1'h0 : _0146_;
  assign _0149_ = _0572_ ? (* src = "CanBsp.scala:368.35|CanBsp.scala:369.14" *) 1'h0 : _0148_;
  assign _0151_ = _0591_ ? (* src = "CanBsp.scala:374.61|CanBsp.scala:375.11" *) 1'h0 : _0150_;
  assign _0154_ = _0614_ ? (* src = "CanBsp.scala:380.67|CanBsp.scala:381.13" *) 1'h0 : _0153_;
  assign _0155_ = _0646_ ? (* src = "CanBsp.scala:386.56|CanBsp.scala:387.8|CanBsp.scala:108.26" *) _0985_ : id;
  assign _0156_ = _0669_ ? (* src = "CanBsp.scala:390.47|CanBsp.scala:391.10|CanBsp.scala:127.28" *) io_sampledBit : rtr1;
  assign _0157_ = _0693_ ? (* src = "CanBsp.scala:394.47|CanBsp.scala:395.10|CanBsp.scala:129.28" *) io_sampledBit : rtr2;
  assign _0158_ = _0696_ ? (* src = "CanBsp.scala:398.46|CanBsp.scala:399.9|CanBsp.scala:128.27" *) io_sampledBit : ide;
  assign _0159_ = _0698_ ? (* src = "CanBsp.scala:402.46|CanBsp.scala:403.13|CanBsp.scala:107.31" *) _0848_ : dataLen;
  assign _0160_ = _0700_ ? (* src = "CanBsp.scala:406.47|CanBsp.scala:407.13|CanBsp.scala:131.31" *) _1374_ : tmpData;
  assign headerLen = io_extendedMode ? (* src = "CanBsp.scala:241.29" *) _0983_ : 3'h2;
  assign _0161_ = _0705_ ? (* src = "CanBsp.scala:418.43|CanBsp.scala:419.13|CanBsp.scala:138.31" *) 3'h0 : byteCnt;
  assign _0163_ = writeDataToTmpFifo ? (* src = "CanBsp.scala:416.28|CanBsp.scala:417.13" *) _0808_ : _0161_;
  assign _0164_ = _0707_ ? (* src = "CanBsp.scala:426.46|CanBsp.scala:427.11|CanBsp.scala:130.29" *) _0812_ : crcIn;
  assign _0165_ = _0719_ ? (* src = "CanBsp.scala:432.44|CanBsp.scala:433.12|CanBsp.scala:106.30" *) _0757_ : bitCnt;
  assign _0166_ = _0717_ ? (* src = "CanBsp.scala:430.132|CanBsp.scala:431.12" *) 6'h00 : _0165_;
  assign _0167_ = rxEof ? (* src = "CanBsp.scala:438.23|CanBsp.scala:439.14|CanBsp.scala:141.30" *) _0852_ : eofCnt;
  assign _0169_ = _0591_ ? (* src = "CanBsp.scala:436.63|CanBsp.scala:437.14" *) 3'h0 : _0167_;
  assign _0170_ = io_samplePoint ? (* src = "CanBsp.scala:435.24|CanBsp.scala:141.30" *) _0169_ : eofCnt;
  assign _0171_ = bitDeStuffReset ? (* src = "CanBsp.scala:445.31|CanBsp.scala:446.19|CanBsp.scala:139.37" *) 1'h0 : bitStuffCntEn;
  assign _0173_ = _1370_ ? (* src = "CanBsp.scala:454.50|CanBsp.scala:455.19|CanBsp.scala:457.19" *) _0800_ : 3'h1;
  assign _1044_ = _1045_ ? (* src = "CanBsp.scala:243.61" *) _1043_ : 4'h7;
  assign _0174_ = bitDeStuff ? (* src = "CanBsp.scala:452.31|CanBsp.scala:453.19" *) 3'h1 : _0173_;
  assign _0175_ = _1368_ ? (* src = "CanBsp.scala:451.46|CanBsp.scala:109.35" *) _0174_ : bitStuffCnt;
  assign _0176_ = bitDeStuffReset ? (* src = "CanBsp.scala:449.25|CanBsp.scala:450.17" *) 3'h1 : _0175_;
  assign _0177_ = _0722_ ? (* src = "CanBsp.scala:466.31|CanBsp.scala:467.21|CanBsp.scala:469.21" *) _0798_ : 3'h1;
  assign _0178_ = bitDeStuffTx ? (* src = "CanBsp.scala:464.33|CanBsp.scala:465.21" *) 3'h1 : _0177_;
  assign _0180_ = _0721_ ? (* src = "CanBsp.scala:463.40|CanBsp.scala:110.37" *) _0178_ : bitStuffCntTx;
  assign _0181_ = _0720_ ? (* src = "CanBsp.scala:461.40|CanBsp.scala:462.19" *) 3'h1 : _0180_;
  assign _0183_ = goRxCrc ? (* src = "CanBsp.scala:473.22|CanBsp.scala:474.15" *) 1'h0 : _0182_;
  assign _0184_ = goRxAck ? (* src = "CanBsp.scala:481.23|CanBsp.scala:482.12|CanBsp.scala:153.30" *) _0810_ : crcErr;
  assign _0185_ = _0724_ ? (* src = "CanBsp.scala:479.40|CanBsp.scala:480.12" *) 1'h0 : _0184_;
  assign limitedDataLenSubOne = remoteRq ? (* src = "CanBsp.scala:243.40" *) 4'hf : _1044_;
  assign _0187_ = _0725_ ? (* src = "CanBsp.scala:485.61|CanBsp.scala:486.19" *) 1'h0 : _0186_;
  assign _0189_ = _0725_ ? (* src = "CanBsp.scala:491.61|CanBsp.scala:492.19" *) 1'h0 : _0188_;
  assign _0192_ = _0726_ ? (* src = "CanBsp.scala:497.40|CanBsp.scala:498.18" *) 1'h0 : _0191_;
  assign _0194_ = _0731_ ? (* src = "CanBsp.scala:503.38|CanBsp.scala:504.18" *) 1'h0 : _0193_;
  assign _0196_ = _0725_ ? (* src = "CanBsp.scala:509.61|CanBsp.scala:510.21" *) 1'h0 : _0195_;
  assign _0198_ = _0725_ ? (* src = "CanBsp.scala:515.61|CanBsp.scala:516.20" *) 1'h0 : _0197_;
  assign _0200_ = resetWrFifo ? (* src = "CanBsp.scala:545.21|CanBsp.scala:546.12" *) 1'h0 : _0199_;
  assign _0202_ = _0739_ ? (* src = "CanBsp.scala:553.38|CanBsp.scala:554.15|CanBsp.scala:161.33" *) _0982_ : { 1'h0, headerCnt };
  assign _0203_ = resetWrFifo ? (* src = "CanBsp.scala:551.21|CanBsp.scala:552.15" *) 4'h0 : _0202_;
  assign _0204_ = wrFifo ? (* src = "CanBsp.scala:559.22|CanBsp.scala:560.13|CanBsp.scala:160.31" *) _0813_ : { 1'h0, dataCnt };
  assign limitedTxCntExt = _1046_ ? (* src = "CanBsp.scala:271.35" *) 6'h3f : _1050_;
  assign _0205_ = resetWrFifo ? (* src = "CanBsp.scala:557.21|CanBsp.scala:558.13" *) 5'h00 : _0204_;
  assign _0833_ = _0832_ ? (* src = "Lookup.scala:33.37" *) _0836_ : tmpFifo_dataForFifo_MPORT_data;
  assign _0834_ = _0831_ ? (* src = "Lookup.scala:33.37" *) _0843_ : _0833_;
  assign _0835_ = _0830_ ? (* src = "Lookup.scala:33.37" *) _0844_ : _0834_;
  assign _0837_ = _0829_ ? (* src = "Lookup.scala:33.37" *) _0845_ : _0835_;
  assign _0838_ = _0828_ ? (* src = "Lookup.scala:33.37" *) _0847_ : _0837_;
  assign _0839_ = _0827_ ? (* src = "Lookup.scala:33.37" *) _0816_ : _0838_;
  assign _0840_ = _0826_ ? (* src = "Lookup.scala:33.37" *) _0817_ : _0839_;
  assign _0841_ = _0825_ ? (* src = "Lookup.scala:33.37" *) _0819_ : _0840_;
  assign _0842_ = _0824_ ? (* src = "Lookup.scala:33.37" *) _0817_ : _0841_;
  assign limitedTxCntStd = _1051_ ? (* src = "CanBsp.scala:272.35" *) 6'h3f : _1055_;
  assign _0207_ = _0741_ ? (* src = "CanBsp.scala:590.64|CanBsp.scala:591.16" *) 1'h0 : _0206_;
  assign _0208_ = _0547_ ? (* src = "CanBsp.scala:598.59|CanBsp.scala:599.15|CanBsp.scala:145.33" *) _0909_ : errorCnt1;
  assign _0209_ = _0743_ ? (* src = "CanBsp.scala:596.64|CanBsp.scala:597.15" *) 3'h0 : _0208_;
  assign _0211_ = _0743_ ? (* src = "CanBsp.scala:602.64|CanBsp.scala:603.26" *) 1'h0 : _0210_;
  assign _0214_ = _0743_ ? (* src = "CanBsp.scala:608.64|CanBsp.scala:609.21" *) 1'h0 : _0213_;
  assign _0215_ = _0551_ ? (* src = "CanBsp.scala:616.44|CanBsp.scala:617.15|CanBsp.scala:146.33" *) _0911_ : errorCnt2;
  assign _0216_ = _0743_ ? (* src = "CanBsp.scala:614.64|CanBsp.scala:615.15" *) 3'h0 : _0215_;
  assign _0217_ = _0556_ ? (* src = "CanBsp.scala:622.95|CanBsp.scala:623.24|CanBsp.scala:147.42" *) _0850_ : delayedDominantCnt;
  assign _0218_ = _0554_ ? (* src = "CanBsp.scala:620.85|CanBsp.scala:621.24" *) 3'h0 : _0217_;
  assign _0219_ = _0562_ ? (* src = "CanBsp.scala:629.78|CanBsp.scala:630.18|CanBsp.scala:632.18" *) _1065_ : 3'h1;
  assign _0001_ = _0544_ ? (* src = "CanBsp.scala:290.35|CanBsp.scala:291.12" *) 1'h0 : _0000_;
  assign _0220_ = _0560_ ? (* src = "CanBsp.scala:628.51|CanBsp.scala:142.34" *) _0219_ : passiveCnt;
  assign _0221_ = _0558_ ? (* src = "CanBsp.scala:626.82|CanBsp.scala:627.16" *) 3'h1 : _0220_;
  assign _0222_ = io_samplePoint ? (* src = "CanBsp.scala:638.30|CanBsp.scala:639.21|CanBsp.scala:183.39" *) 1'h0 : firstCompareBit;
  assign _0005_ = _0563_ ? (* src = "CanBsp.scala:642.46|CanBsp.scala:643.19" *) 1'h0 : _0004_;
  assign _0006_ = _0566_ ? (* src = "CanBsp.scala:650.67|CanBsp.scala:651.18|CanBsp.scala:151.36" *) _1059_ : overloadCnt1;
  assign _0007_ = _0564_ ? (* src = "CanBsp.scala:648.67|CanBsp.scala:649.18" *) 3'h0 : _0006_;
  assign _0009_ = _0564_ ? (* src = "CanBsp.scala:654.67|CanBsp.scala:655.24" *) 1'h0 : _0008_;
  assign _0010_ = _0570_ ? (* src = "CanBsp.scala:662.46|CanBsp.scala:663.18|CanBsp.scala:152.36" *) _1061_ : overloadCnt2;
  assign _0011_ = _0564_ ? (* src = "CanBsp.scala:660.67|CanBsp.scala:661.18" *) 3'h0 : _0010_;
  assign _0013_ = _0573_ ? (* src = "CanBsp.scala:682.29|CanBsp.scala:690.19" *) io_nodeErrorPassive : 1'h1;
  assign _0152_ = _0545_ ? (* src = "CanBsp.scala:296.36|CanBsp.scala:297.11" *) 1'h0 : _0103_;
  assign _0014_ = _0575_ ? (* src = "CanBsp.scala:693.33|CanBsp.scala:694.19|CanBsp.scala:696.19" *) 1'h0 : 1'h1;
  assign _1387_ = _1352_ ? (* src = "CanBsp.scala:722.19" *) _1384_ : _1386_;
  assign _1379_ = _1352_ ? (* src = "CanBsp.scala:728.19" *) _1376_ : _1378_;
  assign _0025_ = rxCrc ? (* src = "CanBsp.scala:723.23|CanBsp.scala:724.13" *) _1389_ : _0024_;
  assign _0026_ = rxData ? (* src = "CanBsp.scala:721.18|CanBsp.scala:722.13" *) _1387_ : _0025_;
  assign _0028_ = rxCrc ? (* src = "CanBsp.scala:733.23|CanBsp.scala:734.13" *) _1389_ : _0027_;
  assign _0030_ = rxData ? (* src = "CanBsp.scala:731.18|CanBsp.scala:732.13" *) _1381_ : _0028_;
  assign txBit = io_extendedMode ? (* src = "CanBsp.scala:720.25" *) _0026_ : _0030_;
  assign _0015_ = io_sendAck ? (* src = "CanBsp.scala:701.30|CanBsp.scala:702.17|CanBsp.scala:704.17" *) 1'h0 : 1'h1;
  assign _0016_ = _0576_ ? (* src = "CanBsp.scala:699.39|CanBsp.scala:700.19" *) _1032_ : _0015_;
  assign _0791_ = io_tx != io_sampledBit;
  assign _0810_ = crcIn != calculatedCrc;
  assign errorCaptureCodeDirection = ~ io_transmitting;
  assign _0970_ = ~ io_nodeBusOff;
  assign _0965_ = ~ io_sampledBit;
  assign _0955_ = ~ _0962_;
  assign _0748_ = ~ io_selfTestMode;
  assign _0793_ = ~ bitErrExc1;
  assign _0795_ = ~ bitErrExc2;
  assign _0780_ = ~ bitErrExc3;
  assign _0769_ = ~ enableErrorCnt2;
  assign _0773_ = ~ enableOverloadCnt2;
  assign _0782_ = ~ bitErrExc4;
  assign _0784_ = ~ bitErrExc5;
  assign _0786_ = ~ bitErrExc6;
  assign _0974_ = ~ bitDeStuff;
  assign _0788_ = ~ io_resetMode;
  assign _1021_ = ~ err;
  assign _0912_ = ~ io_nodeErrorPassive;
  assign _1324_ = ~ bitDeStuffTx;
  assign _1331_ = ~ rxData;
  assign _1326_ = ~ _1352_;
  assign _1332_ = ~ io_extendedMode;
  assign _1027_ = ~ nodeBusOffQ;
  assign _1035_ = ~ errorFrameEnded;
  assign _1037_ = ~ overloadFrameEnded;
  assign _1319_ = ~ ide;
  assign _1039_ = ~ arbitrationLost;
  assign _1030_ = ~ txQ;
  assign _1398_ = ~ goEarlyTxLatched;
  assign _1023_ = ~ arbitrationLostQ;
  assign _1025_ = ~ arbitrationBlocked;
  assign _0626_ = ~ crcErr;
  assign _0633_ = ~ rule5;
  assign _0635_ = ~ errorFlagOverLatched;
  assign _0652_ = ~ _0733_;
  assign _0659_ = ~ _0658_;
  assign _0759_ = ~ io_goErrorFrame;
  assign _1014_ = ~ io_rxIdle;
  assign _1017_ = ~ waitingForBusFree;
  assign _1026_ = ~ errorCaptureCodeBlocked;
  assign io_nodeErrorActive = ~ _1012_;
  assign io_busOffOn = ~ io_nodeBusOff;
  assign _0938_ = ~ io_listenOnlyMode;
  assign _0941_ = ~ io_txState;
  assign _0943_ = ~ suspend;
  assign _0927_ = ~ io_transmitter;
  assign _0957_ = ~ remoteRq;
  assign _0225_ = reset | _0021_;
  assign _0448_ = reset | _0086_;
  assign goRxIdle = _0969_ | _0971_;
  assign _1072_ = _1068_ | _1071_;
  assign _0708_ = goRxRtr2 | io_goErrorFrame;
  assign _0201_ = goRxId2 | rxId2;
  assign _0718_ = goRxR1 | io_goErrorFrame;
  assign _0002_ = goRxRtr2 | rxRtr2;
  assign _0723_ = goRxR0 | io_goErrorFrame;
  assign _0019_ = goRxR1 | rxR1;
  assign _0729_ = goRxDlc | io_goErrorFrame;
  assign _0039_ = goRxR0 | rxR0;
  assign _0735_ = goRxData | goRxCrc;
  assign _0546_ = _0735_ | io_goErrorFrame;
  assign _1078_ = _1074_ | _1077_;
  assign _0061_ = goRxDlc | rxDlc;
  assign _0550_ = goRxCrc | io_goErrorFrame;
  assign _0083_ = goRxData | rxData;
  assign _0557_ = goRxCrcLim | io_goErrorFrame;
  assign _0104_ = goRxCrc | rxCrc;
  assign _0126_ = goRxCrcLim | rxCrcLim;
  assign _0569_ = goRxAckLim | io_goErrorFrame;
  assign _0146_ = goRxAck | rxAck;
  assign _0572_ = goRxEof | io_goErrorFrame;
  assign _0148_ = goRxAckLim | rxAckLim;
  assign _0935_ = _0933_ | _0934_;
  assign _0582_ = io_goRxInter | io_goErrorFrame;
  assign _0591_ = _0582_ | io_goOverloadFrame;
  assign _0150_ = goRxEof | rxEof;
  assign _0600_ = goRxIdle | goRxId1;
  assign _0608_ = _0600_ | io_goOverloadFrame;
  assign _0614_ = _0608_ | io_goErrorFrame;
  assign _0153_ = io_goRxInter | rxInter;
  assign _0621_ = rxId1 | rxId2;
  assign _0709_ = goRxId1 | goRxId2;
  assign _0710_ = _0709_ | goRxDlc;
  assign _0929_ = _0935_ | _0928_;
  assign _0711_ = _0710_ | goRxData;
  assign _0712_ = _0711_ | goRxCrc;
  assign _0713_ = _0712_ | goRxAck;
  assign _0714_ = _0713_ | goRxEof;
  assign _0715_ = _0714_ | io_goRxInter;
  assign _0716_ = _0715_ | io_goErrorFrame;
  assign _0717_ = _0716_ | io_goOverloadFrame;
  assign _0172_ = bitDeStuffSet | _0171_;
  assign _0720_ = io_resetMode | bitDeStuffReset;
  assign _0182_ = goCrcEnable | crcEnable;
  assign _0932_ = _0929_ | _0931_;
  assign _0724_ = io_resetMode | errorFrameEnded;
  assign _0725_ = _0724_ | io_goOverloadFrame;
  assign _0186_ = ackErr | ackErrLatched;
  assign _0188_ = bitErr | bitErrLatched;
  assign _0726_ = io_goErrorFrame | rule3Exc1_1;
  assign _0191_ = _0730_ | rule3Exc1_1;
  assign _0731_ = errorFlagOver | rule3Exc1_1;
  assign _0193_ = _0733_ | rule3Exc1_0;
  assign _0195_ = stuffErr | stuffErrLatched;
  assign _0197_ = formErr | formErrLatched;
  assign _0963_ = io_sampledBit | _0962_;
  assign _0737_ = _0941_ | io_selfRxRequest;
  assign _0199_ = _0738_ | wrFifo;
  assign _0740_ = io_setResetMode | errorFrameEnded;
  assign _0741_ = _0740_ | io_goOverloadFrame;
  assign _0206_ = io_goErrorFrame | errorFrame;
  assign _0742_ = errorFrameEnded | io_goErrorFrame;
  assign _0743_ = _0742_ | io_goOverloadFrame;
  assign _0210_ = errorFlagOver | errorFlagOverLatched;
  assign _0213_ = _0549_ | enableErrorCnt2;
  assign _0552_ = enableErrorCnt2 | io_goErrorFrame;
  assign _0950_ = _0956_ | remoteRq;
  assign _0553_ = _0552_ | enableOverloadCnt2;
  assign _0554_ = _0553_ | io_goOverloadFrame;
  assign _0555_ = _0767_ | _0771_;
  assign _0558_ = _0743_ | firstCompareBit;
  assign _0003_ = io_goErrorFrame | _0222_;
  assign _0563_ = overloadFrameEnded | io_goErrorFrame;
  assign _0004_ = io_goOverloadFrame | overloadFrame;
  assign _0564_ = _0563_ | io_goOverloadFrame;
  assign _0008_ = _0568_ | enableOverloadCnt2;
  assign _0571_ = io_resetMode | io_nodeBusOff;
  assign _0953_ = _0951_ | _0952_;
  assign _0574_ = io_goOverloadFrame | io_overloadFrame;
  assign _0576_ = io_goTx | io_txState;
  assign _0024_ = finishMsg | _1379_;
  assign _0027_ = finishMsg | _1383_;
  assign _1032_ = _1029_ | _1031_;
  assign _0021_ = io_resetMode | _0020_;
  assign _0577_ = io_txState | io_goTx;
  assign _0580_ = goEarlyTx | _0579_;
  assign _0581_ = io_txSuccessful | io_resetMode;
  assign _0584_ = _0581_ | _0583_;
  assign _1007_ = _1006_ | errorFrameEnded;
  assign _0587_ = _0584_ | _0586_;
  assign _0033_ = _0588_ | needToTx;
  assign _1009_ = _0943_ | _1008_;
  assign _1011_ = goEarlyTx | io_rxIdle;
  assign _0589_ = io_resetMode | io_txPoint;
  assign _0035_ = goEarlyTx | goEarlyTxLatched;
  assign _0590_ = io_resetMode | io_goRxInter;
  assign _0592_ = _0590_ | errorFrame;
  assign _0593_ = _0592_ | arbitrationLost;
  assign _0037_ = io_goTx | txState;
  assign resetWrFifo = _1323_ | io_resetMode;
  assign _0594_ = io_resetMode | goRxIdle;
  assign _0596_ = _0594_ | _0595_;
  assign _0041_ = io_goTx | _0040_;
  assign _0597_ = io_goErrorFrame | io_goOverloadFrame;
  assign _0598_ = _0597_ | io_goTx;
  assign _0599_ = _0598_ | io_sendAck;
  assign _0602_ = _0594_ | _0601_;
  assign _0604_ = _0602_ | _0603_;
  assign _0043_ = _0599_ | _0042_;
  assign _0605_ = io_resetMode | _1008_;
  assign _0967_ = io_rxIdle | lastBitOfInter;
  assign _0853_ = formErr | stuffErr;
  assign _0044_ = _0607_ | suspend;
  assign _0046_ = _0610_ | suspendCntEn;
  assign _0612_ = _0600_ | errorFrame;
  assign _0615_ = _0612_ | io_resetMode;
  assign _0051_ = goRxCrcLim | finishMsg;
  assign _0616_ = goRxIdle | errorFrameEnded;
  assign _0053_ = _0620_ | arbitrationLost;
  assign _0059_ = io_setArbitrationLostIrq | arbitrationBlocked;
  assign _0623_ = _0927_ | arbitrationLost;
  assign _0641_ = _0639_ | _0640_;
  assign _0778_ = io_txState | errorFrame;
  assign _0644_ = _0641_ | _0643_;
  assign _0647_ = io_txSuccessful | busFree;
  assign _0650_ = _0643_ | _0640_;
  assign _0661_ = _0650_ | _0660_;
  assign _0663_ = _0661_ | _0662_;
  assign _0670_ = _0667_ | _0668_;
  assign _0672_ = _0742_ | _0671_;
  assign _0076_ = _0674_ | nodeErrorPassive;
  assign _1012_ = io_nodeErrorPassive | io_nodeBusOff;
  assign _0682_ = _0679_ | _0681_;
  assign _0779_ = _0778_ | io_overloadFrame;
  assign _0686_ = _0683_ | _0685_;
  assign _0078_ = _0686_ | nodeBusOff;
  assign _0691_ = _0671_ | _0690_;
  assign _0084_ = _0691_ | _0082_;
  assign _0085_ = _0690_ | waitingForBusFree;
  assign _0860_ = rxCrcLim | rxAck;
  assign _0861_ = _0860_ | rxAckLim;
  assign _0872_ = _0861_ | rxEof;
  assign _0882_ = _0872_ | io_rxInter;
  assign _0892_ = _0882_ | errorFrame;
  assign _0789_ = _0779_ | rxAck;
  assign _0902_ = _0892_ | io_overloadFrame;
  assign _0905_ = _0904_ | rxRtr2;
  assign _0906_ = _0905_ | rxR1;
  assign _0862_ = _0906_ | rxR0;
  assign _0863_ = _0862_ | rxDlc;
  assign _0864_ = _0863_ | rxData;
  assign _0865_ = _0864_ | rxCrc;
  assign _0866_ = _0865_ | rxCrcLim;
  assign _0867_ = _0866_ | rxAck;
  assign _0868_ = _0867_ | rxAckLim;
  assign _0751_ = rxId1 | rxRtr1;
  assign _0869_ = _0868_ | rxEof;
  assign _0870_ = _0869_ | io_overloadFrame;
  assign _0874_ = _0873_ | rxRtr1;
  assign _0875_ = _0874_ | rxIde;
  assign _0876_ = _0875_ | rxId2;
  assign _0877_ = _0876_ | rxRtr2;
  assign _0878_ = _0877_ | rxR1;
  assign _0879_ = _0878_ | _0765_;
  assign _0880_ = _0879_ | io_overloadFrame;
  assign _0881_ = io_rxIdle | rxId1;
  assign _0752_ = _0751_ | rxIde;
  assign _0883_ = _0881_ | rxId2;
  assign _0884_ = _0883_ | rxDlc;
  assign _0885_ = _0884_ | rxData;
  assign _0886_ = _0885_ | rxAckLim;
  assign _0887_ = _0886_ | rxEof;
  assign _0888_ = _0887_ | io_rxInter;
  assign _0889_ = _0888_ | _0765_;
  assign _0890_ = io_rxIdle | rxIde;
  assign _0894_ = _0890_ | _0893_;
  assign _0895_ = _0894_ | rxR1;
  assign _0753_ = _0752_ | rxId2;
  assign _0896_ = _0895_ | rxR0;
  assign _0897_ = _0896_ | rxDlc;
  assign _0898_ = _0897_ | rxAck;
  assign _0899_ = _0898_ | rxAckLim;
  assign _0901_ = _0899_ | _0900_;
  assign _1016_ = waitingForBusFree | _1015_;
  assign _0091_ = io_setBusErrorIrq | errorCaptureCodeBlocked;
  assign _0988_ = _0986_ | _0987_;
  assign _0991_ = _0989_ | _0990_;
  assign io_goRxInter = _1007_ | overloadFrameEnded;
  assign arbitrationField = _0753_ | rxRtr2;
  assign io_transmitStatus = io_transmitting | _1028_;
  assign io_txNext = _0571_ | _0018_;
  assign io_goOverloadFrame = _0996_ | _0998_;
  assign io_goErrorFrame = _0855_ | _0992_;
  assign _0464_ = io_hardSync | io_goTx;
  assign _0467_ = rtr1 | _1056_;
  assign _0468_ = rtr1 | _1057_;
  assign bitErrExc4 = _0770_ | _0774_;
  assign bitErrExc5 = _0775_ | _0776_;
  assign _0973_ = _0972_ | rxR1;
  assign _0854_ = _0853_ | bitErr;
  assign _0855_ = _0854_ | ackErr;
  assign _0856_ = _0855_ | formErrLatched;
  assign _0857_ = _0856_ | stuffErrLatched;
  assign _0858_ = _0857_ | bitErrLatched;
  assign _0859_ = _0858_ | ackErrLatched;
  assign err = _0859_ | crcErr;
  assign _1306_ = _1228_ | _1299_;
  assign _1151_ = _1117_ | _1144_;
  assign rTxData_0 = _1183_ | _1210_;
  assign remoteRq = _1320_ | _1321_;
  assign _1274_ = _1241_ | _1267_;
  assign _1286_ = _1282_ | _1285_;
  assign rTxData_1 = _1289_ | _1292_;
  assign _1298_ = _1294_ | _1297_;
  assign _1305_ = _1301_ | _1304_;
  assign rTxData_2 = _1308_ | _1311_;
  assign _1317_ = _1313_ | _1316_;
  assign _1102_ = _1098_ | _1101_;
  assign rTxData_3 = _1104_ | _1107_;
  assign _1114_ = _1109_ | _1113_;
  assign goCrcEnable = io_hardSync | io_goTx;
  assign _1121_ = _1116_ | _1120_;
  assign rTxData_4 = _1123_ | _1127_;
  assign _1134_ = _1129_ | _1133_;
  assign _1140_ = _1136_ | _1139_;
  assign rTxData_5 = _1142_ | _1146_;
  assign _1153_ = _1148_ | _1152_;
  assign _1159_ = _1155_ | _1158_;
  assign rTxData_6 = _1161_ | _1165_;
  assign _1171_ = _1167_ | _1170_;
  assign _1178_ = _1173_ | _1177_;
  assign _0758_ = goRxAck | io_goErrorFrame;
  assign rTxData_7 = _1180_ | _1184_;
  assign _1191_ = _1186_ | _1189_;
  assign _1198_ = _1193_ | _1196_;
  assign rTxData_8 = _1200_ | _1203_;
  assign _1209_ = _1205_ | _1208_;
  assign _1216_ = _1212_ | _1215_;
  assign rTxData_9 = _1218_ | _1221_;
  assign _1227_ = _1223_ | _1226_;
  assign _1234_ = _1230_ | _1233_;
  assign rTxData_10 = _1237_ | _1240_;
  assign bitDeStuffReset = _0758_ | io_goOverloadFrame;
  assign _1247_ = _1243_ | _1246_;
  assign _1254_ = _1250_ | _1253_;
  assign rTxData_11 = _1257_ | _1260_;
  assign _1266_ = _1262_ | _1265_;
  assign _1273_ = _1269_ | _1272_;
  assign rTxData_12 = _1276_ | _1279_;
  assign _0918_ = _0914_ | _0917_;
  assign _1360_ = _1357_ | _1359_;
  assign _1330_ = _1355_ | _1329_;
  assign _1335_ = _1330_ | _1334_;
  assign _0945_ = _0943_ | _0944_;
  assign _1341_ = _1335_ | _1340_;
  assign _1346_ = _1341_ | _1345_;
  assign _1348_ = _1346_ | _1347_;
  assign _1349_ = goRxIdle | errorFrame;
  assign _1350_ = _1349_ | io_resetMode;
  assign _1351_ = _1350_ | io_overloadFrame;
  assign rstTxPointer = _1348_ | _1351_;
  assign _1001_ = _1000_ | errorFrameEnded;
  assign _1002_ = _1001_ | overloadFrameEnded;
  assign _0996_ = _1003_ | _0995_;
  assign _1097_ = _1088_ | _1096_;
  assign _0997_ = _0919_ | _1063_;
  assign _0544_ = goRxId1 | io_goErrorFrame;
  assign _0000_ = goRxIdle | rxIdle;
  assign _0545_ = goRxRtr1 | io_goErrorFrame;
  assign _0103_ = goRxId1 | rxId1;
  assign _0613_ = goRxIde | io_goErrorFrame;
  assign _0162_ = goRxRtr1 | rxRtr1;
  assign _0692_ = goRxR0 | goRxId2;
  assign _0701_ = _0692_ | io_goErrorFrame;
  assign _0179_ = goRxIde | rxIde;
  always @(posedge clock)
    firstCompareBit <= _1520_;
  always @(posedge clock)
    errorCaptureCodeBlocked <= _1522_;
  always @(posedge clock)
    errorFlagOverLatched <= _1524_;
  always @(posedge clock)
    suspendCnt <= _1526_;
  always @(posedge clock)
    suspendCntEn <= _1528_;
  always @(posedge clock)
    suspend <= _1530_;
  always @(posedge clock)
    rule3Exc1_1 <= _1532_;
  always @(posedge clock)
    rule3Exc1_0 <= _1534_;
  always @(posedge clock)
    formErrLatched <= _1536_;
  always @(posedge clock)
    stuffErrLatched <= _1538_;
  always @(posedge clock)
    bitErrLatched <= _1540_;
  always @(posedge clock)
    ackErrLatched <= _1542_;
  always @(posedge clock)
    nodeBusOffQ <= _1544_;
  always @(posedge clock)
    busFree <= _1546_;
  always @(posedge clock)
    waitingForBusFree <= _0448_;
  always @(posedge clock)
    busFreeCntEn <= _1548_;
  always @(posedge clock)
    busFreeCnt <= _1550_;
  always @(posedge clock)
    finishMsg <= _1552_;
  always @(posedge clock)
    txPointer <= _1554_;
  always @(posedge clock)
    wrFifo <= _1556_;
  always @(posedge clock)
    headerCnt <= _0145_[2:0];
  always @(posedge clock)
    dataCnt <= _0144_[3:0];
  always @(posedge clock)
    txQ <= _1558_;
  always @(posedge clock)
    arbitrationBlocked <= _1560_;
  always @(posedge clock)
    arbitrationCnt <= _1562_;
  always @(posedge clock)
    arbitrationFieldD <= _1402_;
  always @(posedge clock)
    arbitrationLostQ <= _1404_;
  always @(posedge clock)
    arbitrationLost <= _1406_;
  always @(posedge clock)
    crcErr <= _1408_;
  always @(posedge clock)
    overloadCnt2 <= _1410_;
  always @(posedge clock)
    overloadCnt1 <= _1412_;
  always @(posedge clock)
    enableOverloadCnt2 <= _1414_;
  always @(posedge clock)
    delayedDominantCnt <= _1416_;
  always @(posedge clock)
    errorCnt2 <= _1418_;
  always @(posedge clock)
    errorCnt1 <= _1420_;
  always @(posedge clock)
    enableErrorCnt2 <= _1422_;
  always @(posedge clock)
    errorFrame <= _1424_;
  always @(posedge clock)
    passiveCnt <= _1426_;
  always @(posedge clock)
    eofCnt <= _1428_;
  always @(posedge clock)
    crcEnable <= _1430_;
  always @(posedge clock)
    bitStuffCntEn <= _1432_;
  always @(posedge clock)
    byteCnt <= _1434_;
  always @(posedge clock)
    writeDataToTmpFifo <= _1436_;
  always @(posedge clock)
    tmpData <= _1438_;
  always @(posedge clock)
    crcIn <= _1440_;
  always @(posedge clock)
    rtr2 <= _1442_;
  always @(posedge clock)
    ide <= _1444_;
  always @(posedge clock)
    rtr1 <= _1446_;
  always @(posedge clock)
    goEarlyTxLatched <= _1448_;
  always @(posedge clock)
    rxEof <= _1450_;
  always @(posedge clock)
    rxAckLim <= _1452_;
  always @(posedge clock)
    rxAck <= _1454_;
  always @(posedge clock)
    rxCrcLim <= _1456_;
  always @(posedge clock)
    rxCrc <= _1458_;
  always @(posedge clock)
    rxData <= _1460_;
  always @(posedge clock)
    rxDlc <= _1462_;
  always @(posedge clock)
    rxR1 <= _1464_;
  always @(posedge clock)
    rxR0 <= _1466_;
  always @(posedge clock)
    rxRtr2 <= _1468_;
  always @(posedge clock)
    rxId2 <= _1470_;
  always @(posedge clock)
    rxIde <= _1472_;
  always @(posedge clock)
    rxRtr1 <= _1474_;
  always @(posedge clock)
    rxId1 <= _1476_;
  always @(posedge clock)
    txPointQ <= _1478_;
  always @(posedge clock)
    bitStuffCntTx <= _1480_;
  always @(posedge clock)
    bitStuffCnt <= _1482_;
  always @(posedge clock)
    id <= _1484_;
  always @(posedge clock)
    dataLen <= _1486_;
  always @(posedge clock)
    bitCnt <= _1488_;
  always @(posedge clock)
    resetModeQ <= _1490_;
  always @(posedge clock)
    tx <= _0225_;
  always @(posedge clock)
    nodeErrorPassive <= _1492_;
  always @(posedge clock)
    arbitrationLostCapture <= _1494_;
  always @(posedge clock)
    txErrorCount <= _1496_;
  always @(posedge clock)
    rxErrorCount <= _1498_;
  always @(posedge clock)
    needToTx <= _1500_;
  always @(posedge clock)
    nodeBusOff <= _1502_;
  always @(posedge clock)
    rxInter <= _1504_;
  always @(posedge clock)
    transmitter <= _1506_;
  always @(posedge clock)
    transmitting <= _1508_;
  always @(posedge clock)
    rxIdle <= _1510_;
  always @(posedge clock)
    errorCaptureCode <= _1512_;
  always @(posedge clock)
    overloadFrame <= _1514_;
  always @(posedge clock)
    txStateQ <= _1516_;
  always @(posedge clock)
    txState <= _1518_;
  assign _1402_ = _1403_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:156.41" *) 1'h0 : _0055_;
  assign _1404_ = _1405_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:155.40" *) 1'h0 : arbitrationLost;
  assign _1406_ = _1407_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:154.39" *) 1'h0 : _0054_;
  assign _1408_ = _1409_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:153.30" *) 1'h0 : _0185_;
  assign _1410_ = _1411_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:152.36" *) 3'h0 : _0011_;
  assign _1412_ = _1413_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:151.36" *) 3'h0 : _0007_;
  assign _1414_ = _1415_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:148.42" *) 1'h0 : _0009_;
  assign _1416_ = _1417_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:147.42" *) 3'h0 : _0218_;
  assign _1418_ = _1419_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:146.33" *) 3'h0 : _0216_;
  assign _1420_ = _1421_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:145.33" *) 3'h0 : _0209_;
  assign _1422_ = _1423_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:144.39" *) 1'h0 : _0214_;
  assign _1424_ = _1425_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:143.34" *) 1'h0 : _0207_;
  assign _1426_ = _1427_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:142.34" *) 3'h1 : _0221_;
  assign _1428_ = _1429_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:141.30" *) 3'h0 : _0170_;
  assign _1430_ = _1431_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:140.33" *) 1'h0 : _0183_;
  assign _1432_ = _1433_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:139.37" *) 1'h0 : _0172_;
  assign _1434_ = _1435_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:138.31" *) 3'h0 : _0163_;
  assign _1436_ = _1437_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:137.42" *) 1'h0 : _0704_;
  assign _1438_ = _1439_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:131.31" *) 8'h00 : _0160_;
  assign _1440_ = _1441_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:130.29" *) 15'h0000 : _0164_;
  assign _1442_ = _1443_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:129.28" *) 1'h0 : _0157_;
  assign _1444_ = _1445_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:128.27" *) 1'h0 : _0158_;
  assign _1446_ = _1447_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:127.28" *) 1'h0 : _0156_;
  assign _1448_ = _1449_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:126.40" *) 1'h0 : _0036_;
  assign _1450_ = _1451_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:125.29" *) 1'h0 : _0151_;
  assign _1452_ = _1453_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:124.32" *) 1'h0 : _0149_;
  assign _1454_ = _1455_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:123.29" *) 1'h0 : _0147_;
  assign _1456_ = _1457_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:122.32" *) 1'h0 : _0137_;
  assign _1458_ = _1459_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:121.29" *) 1'h0 : _0115_;
  assign _1460_ = _1461_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:120.30" *) 1'h0 : _0092_;
  assign _1462_ = _1463_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:119.29" *) 1'h0 : _0072_;
  assign _1464_ = _1465_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:118.27" *) 1'h0 : _0029_;
  assign _1466_ = _1467_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:117.28" *) 1'h0 : _0050_;
  assign _1468_ = _1469_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:116.30" *) 1'h0 : _0012_;
  assign _1470_ = _1471_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:115.29" *) 1'h0 : _0212_;
  assign _1472_ = _1473_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:114.29" *) 1'h0 : _0190_;
  assign _1474_ = _1475_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:113.30" *) 1'h0 : _0168_;
  assign _1476_ = _1477_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:112.29" *) 1'h0 : _0152_;
  assign _1478_ = _1479_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:111.32" *) 1'h0 : _1395_;
  assign _1480_ = _1481_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:110.37" *) 3'h1 : _0181_;
  assign _1482_ = _1483_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:109.35" *) 3'h1 : _0176_;
  assign _1484_ = _1485_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:108.26" *) 29'h00000000 : _0155_;
  assign _1486_ = _1487_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:107.31" *) 4'h0 : _0159_;
  assign _1488_ = _1489_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:106.30" *) 6'h00 : _0166_;
  assign _1490_ = _1491_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:105.34" *) 1'h0 : io_resetMode;
  assign _1492_ = _1493_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:101.40" *) 1'h0 : _0077_;
  assign _1494_ = _1495_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:99.46" *) 5'h00 : _0058_;
  assign _1496_ = _1497_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:97.36" *) 9'h000 : _0075_;
  assign _1498_ = _1499_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:95.36" *) 9'h000 : _0069_;
  assign _1500_ = _1501_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:93.32" *) 1'h0 : _0034_;
  assign _1502_ = _1503_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:91.34" *) 1'h0 : _0079_;
  assign _1504_ = _1505_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:89.31" *) 1'h0 : _0154_;
  assign _1506_ = _1507_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:87.35" *) 1'h0 : _0041_;
  assign _1508_ = _1509_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:85.36" *) 1'h0 : _0043_;
  assign _1510_ = _1511_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:83.30" *) 1'h0 : _0001_;
  assign _1512_ = _1513_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:81.40" *) 8'h00 : _0088_;
  assign _1514_ = _1515_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:79.37" *) 1'h0 : _0005_;
  assign _1516_ = _1517_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:77.32" *) 1'h0 : _1400_;
  assign _1518_ = _1519_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:75.31" *) 1'h0 : _0038_;
  assign _1520_ = _1521_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:183.39" *) 1'h0 : _0003_;
  assign _1522_ = _1523_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:182.47" *) 1'h0 : _0093_;
  assign _1524_ = _1525_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:180.44" *) 1'h0 : _0211_;
  assign _1526_ = _1527_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:179.34" *) 3'h0 : _0049_;
  assign _1528_ = _1529_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:178.36" *) 1'h0 : _0047_;
  assign _1530_ = _1531_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:177.31" *) 1'h0 : _0045_;
  assign _1532_ = _1533_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:176.38" *) 1'h0 : _0192_;
  assign _1534_ = _1535_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:176.38" *) 1'h0 : _0194_;
  assign _1536_ = _1537_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:175.38" *) 1'h0 : _0198_;
  assign _1538_ = _1539_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:174.39" *) 1'h0 : _0196_;
  assign _1540_ = _1541_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:173.37" *) 1'h0 : _0189_;
  assign _1542_ = _1543_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:172.37" *) 1'h0 : _0187_;
  assign _1544_ = _1545_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:171.35" *) 1'h0 : nodeBusOff;
  assign _1546_ = _1547_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:170.31" *) 1'h0 : _0806_;
  assign _1548_ = _1549_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:168.36" *) 1'h0 : _0084_;
  assign _1550_ = _1551_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:167.34" *) 4'h0 : _0081_;
  assign _1552_ = _1553_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:166.33" *) 1'h0 : _0052_;
  assign _1554_ = _1555_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:164.33" *) 6'h00 : _0032_;
  assign _1556_ = _1557_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:162.30" *) 1'h0 : _0200_;
  assign _1558_ = _1559_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:159.27" *) 1'h0 : _0023_;
  assign _1560_ = _1561_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:158.42" *) 1'h0 : _0060_;
  assign _1562_ = _1563_ ? (* full_case = 32'd1 *) (* src = "CanBsp.scala:157.38" *) 5'h00 : _0057_;
  assign _0919_ = & errorCnt2;
  assign _0767_ = & errorCnt1;
  assign _0703_ = & _0702_;
  assign _0962_ = | _0961_;
  assign _1013_ = | _1040_;
  assign _1375_ = extendedChainDataExt >> txPointer;
  assign _1385_ = extendedChainDataStd >> txPointer;
  assign _1388_ = rCalculatedCrc >> txPointer;
  assign _1390_ = extendedChainExt >> txPointer;
  assign _1377_ = extendedChainStd >> txPointer;
  assign _1380_ = basicChainData >> txPointer;
  assign _1382_ = basicChain >> txPointer;
  assign _0762_ = { 1'h0, _0761_ } - 7'h01;
  assign _1042_ = { 1'h0, dataLen } - 5'h01;
  assign _1049_ = { 1'h0, _1048_ } - 7'h01;
  assign _1054_ = { 1'h0, _1053_ } - 7'h01;
  assign _0815_ = { 1'h0, dataCnt } - { 1'h0, _0814_ };
  assign _1362_ = { 1'h0, io_rxErrorCount } - 10'h001;
  assign _1391_ = { 1'h0, txErrorCount } - 10'h001;
  (* module_not_derived = 32'd1 *)
  (* src = "CanBsp.scala:526.31" *)
  CanAcf canAcf (
    .clock(clock),
    .io_acceptanceCode_0(io_acceptanceCode_0),
    .io_acceptanceCode_1(io_acceptanceCode_1),
    .io_acceptanceCode_2(io_acceptanceCode_2),
    .io_acceptanceCode_3(io_acceptanceCode_3),
    .io_acceptanceFilterMode(io_acceptanceFilterMode),
    .io_acceptanceMask_0(io_acceptanceMask_0),
    .io_acceptanceMask_1(io_acceptanceMask_1),
    .io_acceptanceMask_2(io_acceptanceMask_2),
    .io_acceptanceMask_3(io_acceptanceMask_3),
    .io_data0(tmpFifo_canAcf_io_data0_MPORT_data),
    .io_data1(tmpFifo_canAcf_io_data1_MPORT_data),
    .io_extendedMode(io_extendedMode),
    .io_goErrorFrame(io_goErrorFrame),
    .io_goRxCrcLim(_0466_),
    .io_goRxInter(io_goRxInter),
    .io_id(id),
    .io_idOk(canAcf_io_idOk),
    .io_ide(ide),
    .io_noByte0(_0467_),
    .io_noByte1(_0468_),
    .io_resetMode(io_resetMode),
    .io_rtr1(rtr1),
    .io_rtr2(rtr2),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanBsp.scala:521.72" *)
  CanCrc canCrcRx (
    .clock(clock),
    .io_crc(canCrcRx_io_crc),
    .io_data(io_sampledBit),
    .io_enable(_0465_),
    .reset(_0464_)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanBsp.scala:577.33" *)
  CanFifo canFifo (
    .clock(clock),
    .io_addr(io_addr[5:0]),
    .io_dataIn(_0224_),
    .io_dataOut(canFifo_io_dataOut),
    .io_extendedMode(io_extendedMode),
    .io_infoCnt(canFifo_io_infoCnt),
    .io_infoEmpty(canFifo_io_infoEmpty),
    .io_overrun(canFifo_io_overrun),
    .io_releaseBuffer(io_releaseBuffer),
    .io_resetMode(io_resetMode),
    .io_wr(wrFifo),
    .reset(reset)
  );
  assign _1040_ = bitCnt[1:0];
  assign _0977_ = bitCnt[3:0];
  assign _0980_ = bitCnt[4:0];
  assign calculatedCrc = canCrcRx_io_crc;
  assign _1066_ = calculatedCrc[7:0];
  assign _1079_ = _1066_[7:4];
  assign _0094_ = { 4'h0, _1079_ };
  assign _1094_ = _1066_[3:0];
  assign _1095_ = { _1094_, 4'h0 };
  assign _1067_ = _1097_[7:2];
  assign _0095_ = { 2'h0, _1067_ };
  assign _1069_ = _1097_[5:0];
  assign _1070_ = { _1069_, 2'h0 };
  assign _1073_ = _1072_[7:1];
  assign _0096_ = { 1'h0, _1073_ };
  assign _1075_ = _1072_[6:0];
  assign _1076_ = { _1075_, 1'h0 };
  assign _1080_ = calculatedCrc[14:8];
  assign _1081_ = _1080_[3:0];
  assign _1082_ = _1081_[1:0];
  assign _1083_ = _1082_[0];
  assign _1084_ = _1082_[1];
  assign _1085_ = _1081_[3:2];
  assign _1086_ = _1085_[0];
  assign _1087_ = _1085_[1];
  assign _1089_ = _1080_[6:4];
  assign _1090_ = _1089_[1:0];
  assign _1091_ = _1090_[0];
  assign _1092_ = _1090_[1];
  assign _1093_ = _1089_[2];
  assign rCalculatedCrc = { _1078_, _1083_, _1084_, _1086_, _1087_, _1091_, _1092_, _1093_ };
  assign _0760_ = limitedDataLen[2:0];
  assign _0761_ = { _0760_, 3'h0 };
  assign _0763_ = _0762_[5:0];
  assign _0961_ = dataLen[2:0];
  assign _1043_ = _1042_[3:0];
  assign _0097_ = { 1'h0, headerLen };
  assign _0098_ = { 1'h0, dataCnt };
  assign _1164_ = io_txData_0[7:4];
  assign _0099_ = { 4'h0, _1164_ };
  assign _1280_ = io_txData_0[3:0];
  assign _1287_ = { _1280_, 4'h0 };
  assign _1110_ = _1306_[7:2];
  assign _0100_ = { 2'h0, _1110_ };
  assign _1124_ = _1306_[5:0];
  assign _1131_ = { _1124_, 2'h0 };
  assign _1176_ = _1151_[7:1];
  assign _0101_ = { 1'h0, _1176_ };
  assign _1190_ = _1151_[6:0];
  assign _1197_ = { _1190_, 1'h0 };
  assign _1235_ = io_txData_1[7:4];
  assign _0102_ = { 4'h0, _1235_ };
  assign _1248_ = io_txData_1[3:0];
  assign _1255_ = { _1248_, 4'h0 };
  assign _1281_ = _1274_[7:2];
  assign _0105_ = { 2'h0, _1281_ };
  assign _1283_ = _1274_[5:0];
  assign _1284_ = { _1283_, 2'h0 };
  assign _1288_ = _1286_[7:1];
  assign _0106_ = { 1'h0, _1288_ };
  assign _1290_ = _1286_[6:0];
  assign _1291_ = { _1290_, 1'h0 };
  assign _1293_ = io_txData_2[7:4];
  assign _0107_ = { 4'h0, _1293_ };
  assign _1295_ = io_txData_2[3:0];
  assign _1296_ = { _1295_, 4'h0 };
  assign _1300_ = _1298_[7:2];
  assign _0108_ = { 2'h0, _1300_ };
  assign _1302_ = _1298_[5:0];
  assign _1303_ = { _1302_, 2'h0 };
  assign _1307_ = _1305_[7:1];
  assign _0109_ = { 1'h0, _1307_ };
  assign _1309_ = _1305_[6:0];
  assign _1310_ = { _1309_, 1'h0 };
  assign _1312_ = io_txData_3[7:4];
  assign _0110_ = { 4'h0, _1312_ };
  assign _1314_ = io_txData_3[3:0];
  assign _1315_ = { _1314_, 4'h0 };
  assign _1318_ = _1317_[7:2];
  assign _0111_ = { 2'h0, _1318_ };
  assign _1099_ = _1317_[5:0];
  assign _1100_ = { _1099_, 2'h0 };
  assign _1103_ = _1102_[7:1];
  assign _0112_ = { 1'h0, _1103_ };
  assign _1105_ = _1102_[6:0];
  assign _1106_ = { _1105_, 1'h0 };
  assign _1108_ = io_txData_4[7:4];
  assign _0113_ = { 4'h0, _1108_ };
  assign _1111_ = io_txData_4[3:0];
  assign _1112_ = { _1111_, 4'h0 };
  assign _1115_ = _1114_[7:2];
  assign _0114_ = { 2'h0, _1115_ };
  assign _1118_ = _1114_[5:0];
  assign _1119_ = { _1118_, 2'h0 };
  assign _1122_ = _1121_[7:1];
  assign _0116_ = { 1'h0, _1122_ };
  assign _1125_ = _1121_[6:0];
  assign _1126_ = { _1125_, 1'h0 };
  assign _1128_ = io_txData_5[7:4];
  assign _0117_ = { 4'h0, _1128_ };
  assign _1130_ = io_txData_5[3:0];
  assign _1132_ = { _1130_, 4'h0 };
  assign _1135_ = _1134_[7:2];
  assign _0118_ = { 2'h0, _1135_ };
  assign _1137_ = _1134_[5:0];
  assign _1138_ = { _1137_, 2'h0 };
  assign _1141_ = _1140_[7:1];
  assign _0119_ = { 1'h0, _1141_ };
  assign _1143_ = _1140_[6:0];
  assign _1145_ = { _1143_, 1'h0 };
  assign _1147_ = io_txData_6[7:4];
  assign _0120_ = { 4'h0, _1147_ };
  assign _1149_ = io_txData_6[3:0];
  assign _1150_ = { _1149_, 4'h0 };
  assign _1154_ = _1153_[7:2];
  assign _0121_ = { 2'h0, _1154_ };
  assign _1156_ = _1153_[5:0];
  assign _1157_ = { _1156_, 2'h0 };
  assign _1160_ = _1159_[7:1];
  assign _0122_ = { 1'h0, _1160_ };
  assign _1162_ = _1159_[6:0];
  assign _1163_ = { _1162_, 1'h0 };
  assign _1166_ = io_txData_7[7:4];
  assign _0123_ = { 4'h0, _1166_ };
  assign _1168_ = io_txData_7[3:0];
  assign _1169_ = { _1168_, 4'h0 };
  assign _1172_ = _1171_[7:2];
  assign _0124_ = { 2'h0, _1172_ };
  assign _1174_ = _1171_[5:0];
  assign _1175_ = { _1174_, 2'h0 };
  assign _1179_ = _1178_[7:1];
  assign _0125_ = { 1'h0, _1179_ };
  assign _1181_ = _1178_[6:0];
  assign _1182_ = { _1181_, 1'h0 };
  assign _1185_ = io_txData_8[7:4];
  assign _0127_ = { 4'h0, _1185_ };
  assign _1187_ = io_txData_8[3:0];
  assign _1188_ = { _1187_, 4'h0 };
  assign _1192_ = _1191_[7:2];
  assign _0128_ = { 2'h0, _1192_ };
  assign _1194_ = _1191_[5:0];
  assign _1195_ = { _1194_, 2'h0 };
  assign _1199_ = _1198_[7:1];
  assign _0129_ = { 1'h0, _1199_ };
  assign _1201_ = _1198_[6:0];
  assign _1202_ = { _1201_, 1'h0 };
  assign _1204_ = io_txData_9[7:4];
  assign _0130_ = { 4'h0, _1204_ };
  assign _1206_ = io_txData_9[3:0];
  assign _1207_ = { _1206_, 4'h0 };
  assign _1211_ = _1209_[7:2];
  assign _0131_ = { 2'h0, _1211_ };
  assign _1213_ = _1209_[5:0];
  assign _1214_ = { _1213_, 2'h0 };
  assign _1217_ = _1216_[7:1];
  assign _0132_ = { 1'h0, _1217_ };
  assign _1219_ = _1216_[6:0];
  assign _1220_ = { _1219_, 1'h0 };
  assign _1222_ = io_txData_10[7:4];
  assign _0133_ = { 4'h0, _1222_ };
  assign _1224_ = io_txData_10[3:0];
  assign _1225_ = { _1224_, 4'h0 };
  assign _1229_ = _1227_[7:2];
  assign _0134_ = { 2'h0, _1229_ };
  assign _1231_ = _1227_[5:0];
  assign _1232_ = { _1231_, 2'h0 };
  assign _1236_ = _1234_[7:1];
  assign _0135_ = { 1'h0, _1236_ };
  assign _1238_ = _1234_[6:0];
  assign _1239_ = { _1238_, 1'h0 };
  assign _1242_ = io_txData_11[7:4];
  assign _0136_ = { 4'h0, _1242_ };
  assign _1244_ = io_txData_11[3:0];
  assign _1245_ = { _1244_, 4'h0 };
  assign _1249_ = _1247_[7:2];
  assign _0138_ = { 2'h0, _1249_ };
  assign _1251_ = _1247_[5:0];
  assign _1252_ = { _1251_, 2'h0 };
  assign _1256_ = _1254_[7:1];
  assign _0139_ = { 1'h0, _1256_ };
  assign _1258_ = _1254_[6:0];
  assign _1259_ = { _1258_, 1'h0 };
  assign _1261_ = io_txData_12[7:4];
  assign _0140_ = { 4'h0, _1261_ };
  assign _1263_ = io_txData_12[3:0];
  assign _1264_ = { _1263_, 4'h0 };
  assign _1268_ = _1266_[7:2];
  assign _0141_ = { 2'h0, _1268_ };
  assign _1270_ = _1266_[5:0];
  assign _1271_ = { _1270_, 2'h0 };
  assign _1275_ = _1273_[7:1];
  assign _0142_ = { 1'h0, _1275_ };
  assign _1277_ = _1273_[6:0];
  assign _1278_ = { _1277_, 1'h0 };
  assign _0754_ = rTxData_1[7:4];
  assign _0755_ = rTxData_1[3:0];
  assign basicChain = { _0754_, 2'h0, _0755_, rTxData_0, 1'h0 };
  assign basicChainData = { rTxData_9, rTxData_8, rTxData_7, rTxData_6, rTxData_5, rTxData_4, rTxData_3, rTxData_2 };
  assign _0922_ = rTxData_0[7:4];
  assign _0923_ = rTxData_0[1];
  assign _0924_ = rTxData_2[2:0];
  assign extendedChainStd = { _0922_, 2'h0, _0923_, _0924_, rTxData_1, 1'h0 };
  assign _0920_ = rTxData_4[4:0];
  assign _0921_ = rTxData_2[7:3];
  assign extendedChainExt = { _0922_, 2'h0, _0923_, _0920_, rTxData_3, _0921_, 2'h3, _0924_, rTxData_1, 1'h0 };
  assign extendedChainDataStd = { rTxData_10, rTxData_9, rTxData_8, rTxData_7, rTxData_6, rTxData_5, rTxData_4, rTxData_3 };
  assign extendedChainDataExt = { rTxData_12, rTxData_11, rTxData_10, rTxData_9, rTxData_8, rTxData_7, rTxData_6, rTxData_5 };
  assign _1046_ = io_txData_0[3];
  assign _1047_ = io_txData_0[2:0];
  assign _1048_ = { _1047_, 3'h0 };
  assign _1050_ = _1049_[5:0];
  assign _1051_ = io_txData_1[3];
  assign _1052_ = io_txData_1[2:0];
  assign _1053_ = { _1052_, 3'h0 };
  assign _1055_ = _1054_[5:0];
  assign _1352_ = rTxData_0[0];
  assign _0984_ = id[27:0];
  assign _0985_ = { _0984_, io_sampledBit };
  assign _0848_ = { _0961_, io_sampledBit };
  assign _1373_ = tmpData[6:0];
  assign _1374_ = { _1373_, io_sampledBit };
  assign _0702_ = bitCnt[2:0];
  assign _0808_ = _0807_[2:0];
  assign _0811_ = crcIn[13:0];
  assign _0812_ = { _0811_, io_sampledBit };
  assign _0757_ = _0756_[5:0];
  assign _0852_ = _0851_[2:0];
  assign _0800_ = _0799_[2:0];
  assign _0798_ = _0797_[2:0];
  assign idOk = canAcf_io_idOk;
  assign fifoSelector = { storingHeader, io_extendedMode, ide, headerCnt };
  assign _0814_ = { 1'h0, headerLen };
  assign _0823_ = _0815_[3:0];
  assign _0836_ = { 1'h1, rtr2, 2'h0, dataLen };
  assign _0843_ = id[28:21];
  assign _0844_ = id[20:13];
  assign _0845_ = id[12:5];
  assign _0846_ = id[4:0];
  assign _0847_ = { _0846_, 3'h0 };
  assign _0816_ = { 1'h0, rtr1, 2'h0, dataLen };
  assign _0817_ = id[10:3];
  assign _0818_ = id[2:0];
  assign _0819_ = { _0818_, rtr1, 4'h0 };
  assign _0820_ = { _0818_, rtr1, dataLen };
  assign _0909_ = _0908_[2:0];
  assign _0911_ = _0910_[2:0];
  assign _0850_ = _0849_[2:0];
  assign _1065_ = _1064_[2:0];
  assign _1059_ = _1058_[2:0];
  assign _1061_ = _1060_[2:0];
  assign _1384_ = _1375_[0];
  assign _1386_ = _1385_[0];
  assign _1389_ = _1388_[0];
  assign _1376_ = _1390_[0];
  assign _1378_ = _1377_[0];
  assign _1381_ = _1380_[0];
  assign _1383_ = _1382_[0];
  assign _1397_ = _1396_[5:0];
  assign _1372_ = _1371_[2:0];
  assign _0750_ = _0749_[4:0];
  assign _1361_ = { 1'h0, io_dataIn };
  assign _1363_ = _1362_[8:0];
  assign _1365_ = _1364_[8:0];
  assign _1367_ = _1366_[8:0];
  assign _1392_ = _1391_[8:0];
  assign _1394_ = _1393_[8:0];
  assign _0802_ = _0801_[3:0];
  assign _0907_ = { errorCaptureCodeType, errorCaptureCodeDirection, _0902_, _0870_, _0880_, _0889_, _0901_ };
  assign _0143_ = { 1'h0, io_errorWarningLimit };
  assign io_dataOut = canFifo_io_dataOut;
  assign io_txState = txState;
  assign io_txStateQ = txStateQ;
  assign io_overloadFrame = overloadFrame;
  assign io_errorCaptureCode = errorCaptureCode;
  assign io_rxIdle = rxIdle;
  assign io_transmitting = transmitting;
  assign io_transmitter = transmitter;
  assign io_rxInter = rxInter;
  assign io_nodeBusOff = nodeBusOff;
  assign io_rxErrorCount = rxErrorCount;
  assign io_txErrorCount = txErrorCount;
  assign io_needToTx = needToTx;
  assign io_overrun = canFifo_io_overrun;
  assign io_infoEmpty = canFifo_io_infoEmpty;
  assign io_arbitrationLostCapture = arbitrationLostCapture;
  assign io_nodeErrorPassive = nodeErrorPassive;
  assign io_rxMessageCounter = canFifo_io_infoCnt;
  assign io_tx = tx;
  assign \waitingForBusFree$process$CanBsp_69  = _0448_;
  assign \headerCnt$process$CanBsp_63  = _0145_[2:0];
  assign \dataCnt$process$CanBsp_62  = _0144_[3:0];
  assign \tx$process$CanBsp_13  = _0225_;
  assign _1521_ = reset;
  assign \firstCompareBit$process$CanBsp_83  = _1520_;
  assign _1523_ = reset;
  assign \errorCaptureCodeBlocked$process$CanBsp_82  = _1522_;
  assign _1525_ = reset;
  assign \errorFlagOverLatched$process$CanBsp_81  = _1524_;
  assign _1527_ = reset;
  assign \suspendCnt$process$CanBsp_80  = _1526_;
  assign _1529_ = reset;
  assign \suspendCntEn$process$CanBsp_79  = _1528_;
  assign _1531_ = reset;
  assign \suspend$process$CanBsp_78  = _1530_;
  assign _1533_ = reset;
  assign \rule3Exc1_1$process$CanBsp_77  = _1532_;
  assign _1535_ = reset;
  assign \rule3Exc1_0$process$CanBsp_76  = _1534_;
  assign _1537_ = reset;
  assign \formErrLatched$process$CanBsp_75  = _1536_;
  assign _1539_ = reset;
  assign \stuffErrLatched$process$CanBsp_74  = _1538_;
  assign _1541_ = reset;
  assign \bitErrLatched$process$CanBsp_73  = _1540_;
  assign _1543_ = reset;
  assign \ackErrLatched$process$CanBsp_72  = _1542_;
  assign _1545_ = reset;
  assign \nodeBusOffQ$process$CanBsp_71  = _1544_;
  assign _1547_ = reset;
  assign \busFree$process$CanBsp_70  = _1546_;
  assign _1549_ = reset;
  assign \busFreeCntEn$process$CanBsp_68  = _1548_;
  assign _1551_ = reset;
  assign \busFreeCnt$process$CanBsp_67  = _1550_;
  assign _1553_ = reset;
  assign \finishMsg$process$CanBsp_66  = _1552_;
  assign _1555_ = reset;
  assign \txPointer$process$CanBsp_65  = _1554_;
  assign _1557_ = reset;
  assign \wrFifo$process$CanBsp_64  = _1556_;
  assign _1559_ = reset;
  assign \txQ$process$CanBsp_61  = _1558_;
  assign _1561_ = reset;
  assign \arbitrationBlocked$process$CanBsp_60  = _1560_;
  assign _1563_ = reset;
  assign \arbitrationCnt$process$CanBsp_59  = _1562_;
  assign _1403_ = reset;
  assign \arbitrationFieldD$process$CanBsp_58  = _1402_;
  assign _1405_ = reset;
  assign \arbitrationLostQ$process$CanBsp_57  = _1404_;
  assign _1407_ = reset;
  assign \arbitrationLost$process$CanBsp_56  = _1406_;
  assign _1409_ = reset;
  assign \crcErr$process$CanBsp_55  = _1408_;
  assign _1411_ = reset;
  assign \overloadCnt2$process$CanBsp_54  = _1410_;
  assign _1413_ = reset;
  assign \overloadCnt1$process$CanBsp_53  = _1412_;
  assign _1415_ = reset;
  assign \enableOverloadCnt2$process$CanBsp_52  = _1414_;
  assign _1417_ = reset;
  assign \delayedDominantCnt$process$CanBsp_51  = _1416_;
  assign _1419_ = reset;
  assign \errorCnt2$process$CanBsp_50  = _1418_;
  assign _1421_ = reset;
  assign \errorCnt1$process$CanBsp_49  = _1420_;
  assign _1423_ = reset;
  assign \enableErrorCnt2$process$CanBsp_48  = _1422_;
  assign _1425_ = reset;
  assign \errorFrame$process$CanBsp_47  = _1424_;
  assign _1427_ = reset;
  assign \passiveCnt$process$CanBsp_46  = _1426_;
  assign _1429_ = reset;
  assign \eofCnt$process$CanBsp_45  = _1428_;
  assign _1431_ = reset;
  assign \crcEnable$process$CanBsp_44  = _1430_;
  assign _1433_ = reset;
  assign \bitStuffCntEn$process$CanBsp_43  = _1432_;
  assign _1435_ = reset;
  assign \byteCnt$process$CanBsp_42  = _1434_;
  assign _1437_ = reset;
  assign \writeDataToTmpFifo$process$CanBsp_41  = _1436_;
  assign _1439_ = reset;
  assign \tmpData$process$CanBsp_40  = _1438_;
  assign _1441_ = reset;
  assign \crcIn$process$CanBsp_39  = _1440_;
  assign _1443_ = reset;
  assign \rtr2$process$CanBsp_38  = _1442_;
  assign _1445_ = reset;
  assign \ide$process$CanBsp_37  = _1444_;
  assign _1447_ = reset;
  assign \rtr1$process$CanBsp_36  = _1446_;
  assign _1449_ = reset;
  assign \goEarlyTxLatched$process$CanBsp_35  = _1448_;
  assign _1451_ = reset;
  assign \rxEof$process$CanBsp_34  = _1450_;
  assign _1453_ = reset;
  assign \rxAckLim$process$CanBsp_33  = _1452_;
  assign _1455_ = reset;
  assign \rxAck$process$CanBsp_32  = _1454_;
  assign _1457_ = reset;
  assign \rxCrcLim$process$CanBsp_31  = _1456_;
  assign _1459_ = reset;
  assign \rxCrc$process$CanBsp_30  = _1458_;
  assign _1461_ = reset;
  assign \rxData$process$CanBsp_29  = _1460_;
  assign _1463_ = reset;
  assign \rxDlc$process$CanBsp_28  = _1462_;
  assign _1465_ = reset;
  assign \rxR1$process$CanBsp_27  = _1464_;
  assign _1467_ = reset;
  assign \rxR0$process$CanBsp_26  = _1466_;
  assign _1469_ = reset;
  assign \rxRtr2$process$CanBsp_25  = _1468_;
  assign _1471_ = reset;
  assign \rxId2$process$CanBsp_24  = _1470_;
  assign _1473_ = reset;
  assign \rxIde$process$CanBsp_23  = _1472_;
  assign _1475_ = reset;
  assign \rxRtr1$process$CanBsp_22  = _1474_;
  assign _1477_ = reset;
  assign \rxId1$process$CanBsp_21  = _1476_;
  assign _1479_ = reset;
  assign \txPointQ$process$CanBsp_20  = _1478_;
  assign _1481_ = reset;
  assign \bitStuffCntTx$process$CanBsp_19  = _1480_;
  assign _1483_ = reset;
  assign \bitStuffCnt$process$CanBsp_18  = _1482_;
  assign _1485_ = reset;
  assign \id$process$CanBsp_17  = _1484_;
  assign _1487_ = reset;
  assign \dataLen$process$CanBsp_16  = _1486_;
  assign _1489_ = reset;
  assign \bitCnt$process$CanBsp_15  = _1488_;
  assign _1491_ = reset;
  assign \resetModeQ$process$CanBsp_14  = _1490_;
  assign _1493_ = reset;
  assign \nodeErrorPassive$process$CanBsp_12  = _1492_;
  assign _1495_ = reset;
  assign \arbitrationLostCapture$process$CanBsp_11  = _1494_;
  assign _1497_ = reset;
  assign \txErrorCount$process$CanBsp_10  = _1496_;
  assign _1499_ = reset;
  assign \rxErrorCount$process$CanBsp_9  = _1498_;
  assign _1501_ = reset;
  assign \needToTx$process$CanBsp_8  = _1500_;
  assign _1503_ = reset;
  assign \nodeBusOff$process$CanBsp_7  = _1502_;
  assign _1505_ = reset;
  assign \rxInter$process$CanBsp_6  = _1504_;
  assign _1507_ = reset;
  assign \transmitter$process$CanBsp_5  = _1506_;
  assign _1509_ = reset;
  assign \transmitting$process$CanBsp_4  = _1508_;
  assign _1511_ = reset;
  assign \rxIdle$process$CanBsp_3  = _1510_;
  assign _1513_ = reset;
  assign \errorCaptureCode$process$CanBsp_2  = _1512_;
  assign _1515_ = reset;
  assign \overloadFrame$process$CanBsp_1  = _1514_;
  assign _1517_ = reset;
  assign \txStateQ$process$CanBsp_0  = _1516_;
  assign _1519_ = reset;
  assign \txState$process$CanBsp  = _1518_;
endmodule

(* cells_not_processed =  1  *)
module CanBtl(clock, reset, io_rx, io_tx, io_baudRatePrescaler, io_syncJumpWidth, io_timeSegment1, io_timeSegment2, io_tripleSampling, io_rxIdle, io_rxInter, io_transmitting, io_transmitter, io_goRxInter, io_txNext, io_goOverloadFrame, io_goErrorFrame, io_goTx, io_sendAck, io_nodeErrorPassive, io_samplePoint
, io_sampledBit, io_sampledBitQ, io_txPoint, io_hardSync);
  (* src = "CanBtl.scala:155.46|CanBtl.scala:156.16|CanBtl.scala:158.16" *)
  wire [6:0] _000_;
  (* src = "CanBtl.scala:195.24|CanBtl.scala:197.19|CanBtl.scala:114.37" *)
  wire [5:0] _001_;
  (* src = "CanBtl.scala:192.34|CanBtl.scala:194.19" *)
  wire [5:0] _002_;
  (* src = "CanBtl.scala:203.30|CanBtl.scala:204.11|CanBtl.scala:116.29" *)
  wire [3:0] _003_;
  (* src = "CanBtl.scala:200.94|CanBtl.scala:201.11" *)
  wire [5:0] _004_;
  (* src = "CanBtl.scala:213.31|CanBtl.scala:214.20|CanBtl.scala:216.20" *)
  wire _005_;
  (* src = "CanBtl.scala:212.65|CanBtl.scala:99.34" *)
  wire _006_;
  (* src = "CanBtl.scala:212.65|CanBtl.scala:218.19|CanBtl.scala:95.35" *)
  wire _007_;
  (* src = "CanBtl.scala:212.65|CanBtl.scala:219.19|CanBtl.scala:101.35" *)
  wire _008_;
  (* src = "CanBtl.scala:211.38|CanBtl.scala:99.34" *)
  wire _009_;
  (* src = "CanBtl.scala:211.38|CanBtl.scala:222.17" *)
  wire _010_;
  (* src = "CanBtl.scala:169.22|CanBtl.scala:170.19|CanBtl.scala:124.37" *)
  wire _011_;
  (* src = "CanBtl.scala:211.38|CanBtl.scala:101.35" *)
  wire _012_;
  (* src = "CanBtl.scala:207.25|CanBtl.scala:208.17" *)
  wire _013_;
  (* src = "CanBtl.scala:207.25|CanBtl.scala:209.17" *)
  wire _014_;
  (* src = "CanBtl.scala:207.25|CanBtl.scala:99.34" *)
  wire _015_;
  (* src = "CanBtl.scala:231.26|CanBtl.scala:232.14|CanBtl.scala:128.31" *)
  wire _016_;
  (* src = "CanBtl.scala:228.52|CanBtl.scala:229.14" *)
  wire _017_;
  (* src = "CanBtl.scala:225.94|CanBtl.scala:226.14" *)
  wire _018_;
  (* src = "CanBtl.scala:238.24|CanBtl.scala:239.19|CanBtl.scala:110.35" *)
  wire _019_;
  (* src = "CanBtl.scala:236.18|CanBtl.scala:237.19" *)
  wire _020_;
  (* src = "CanBtl.scala:235.18|CanBtl.scala:110.35" *)
  wire _021_;
  (* src = "CanBtl.scala:167.37|CanBtl.scala:168.19" *)
  wire _022_;
  (* src = "CanBtl.scala:246.84|CanBtl.scala:247.21|CanBtl.scala:112.39" *)
  wire _023_;
  (* src = "CanBtl.scala:243.107|CanBtl.scala:244.21" *)
  wire _024_;
  (* src = "CanBtl.scala:151.77" *)
  wire [3:0] _025_;
  (* src = "CanBtl.scala:151.57" *)
  wire [3:0] _026_;
  (* src = "CanBtl.scala:155.19" *)
  wire [7:0] _027_;
  (* src = "CanBtl.scala:201.32" *)
  wire [4:0] _028_;
  (* src = "CanBtl.scala:114.37|CanBtl.scala:114.37" *)
  wire [5:0] _029_;
  (* src = "CanBtl.scala:116.29|CanBtl.scala:116.29" *)
  wire [5:0] _030_;
  (* src = "CanBtl.scala:173.18|CanBtl.scala:174.10|CanBtl.scala:118.28" *)
  wire _031_;
  (* src = "CanBtl.scala:173.18|CanBtl.scala:175.12|CanBtl.scala:126.30" *)
  wire [1:0] _032_;
  (* src = "CanBtl.scala:181.22|CanBtl.scala:183.10|CanBtl.scala:120.28" *)
  wire _033_;
  (* src = "CanBtl.scala:178.16|CanBtl.scala:180.10" *)
  wire _034_;
  (* src = "CanBtl.scala:188.31|CanBtl.scala:189.10|CanBtl.scala:122.28" *)
  wire _035_;
  (* src = "CanBtl.scala:186.16|CanBtl.scala:187.10" *)
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire [4:0] _040_;
  wire [3:0] _041_;
  wire _042_;
  wire [5:0] _043_;
  wire [5:0] _044_;
  wire [5:0] _045_;
  (* src = "CanBtl.scala:155.38" *)
  wire [8:0] _046_;
  (* src = "CanBtl.scala:155.38" *)
  wire [7:0] _047_;
  (* src = "CanBtl.scala:192.24" *)
  wire _048_;
  (* src = "CanBtl.scala:200.15" *)
  wire _049_;
  (* src = "CanBtl.scala:200.25" *)
  wire _050_;
  (* src = "CanBtl.scala:200.81" *)
  wire _051_;
  (* src = "CanBtl.scala:200.72" *)
  wire _052_;
  (* src = "CanBtl.scala:200.60" *)
  wire _053_;
  (* src = "CanBtl.scala:200.42" *)
  wire _054_;
  (* src = "CanBtl.scala:200.22" *)
  wire _055_;
  (* src = "CanBtl.scala:155.19" *)
  wire _056_;
  (* src = "CanBtl.scala:211.22" *)
  wire _057_;
  (* src = "CanBtl.scala:212.15" *)
  wire _058_;
  (* src = "CanBtl.scala:225.48" *)
  wire _059_;
  (* src = "CanBtl.scala:225.46" *)
  wire _060_;
  (* src = "CanBtl.scala:225.27" *)
  wire _061_;
  (* src = "CanBtl.scala:225.70" *)
  wire _062_;
  (* src = "CanBtl.scala:225.80" *)
  wire _063_;
  (* src = "CanBtl.scala:228.29" *)
  wire _064_;
  (* src = "CanBtl.scala:243.20" *)
  wire _065_;
  (* src = "CanBtl.scala:243.50" *)
  wire _066_;
  (* src = "CanBtl.scala:243.67" *)
  wire _067_;
  (* src = "CanBtl.scala:243.78" *)
  wire _068_;
  (* src = "CanBtl.scala:243.94" *)
  wire _069_;
  (* src = "CanBtl.scala:243.91" *)
  wire _070_;
  (* src = "CanBtl.scala:243.31" *)
  wire _071_;
  (* src = "CanBtl.scala:246.53" *)
  wire _072_;
  (* src = "CanBtl.scala:246.67" *)
  wire _073_;
  (* src = "CanBtl.scala:246.26" *)
  wire _074_;
  (* src = "CanBtl.scala:161.19" *)
  wire _075_;
  (* src = "CanBtl.scala:167.24" *)
  wire _076_;
  (* src = "CanBtl.scala:167.22" *)
  wire _077_;
  (* src = "CanBtl.scala:188.21" *)
  wire _078_;
  (* src = "CanBtl.scala:158.30" *)
  wire [7:0] _079_;
  (* src = "CanBtl.scala:158.30" *)
  wire [6:0] _080_;
  (* src = "CanBtl.scala:201.32" *)
  wire _081_;
  (* src = "CanBtl.scala:201.17" *)
  wire [5:0] _082_;
  (* src = "CanBtl.scala:138.40" *)
  wire _083_;
  (* src = "CanBtl.scala:138.64" *)
  wire _084_;
  (* src = "CanBtl.scala:138.71" *)
  wire _085_;
  (* src = "CanBtl.scala:138.54" *)
  wire _086_;
  (* src = "CanBtl.scala:138.102" *)
  wire _087_;
  (* src = "CanBtl.scala:138.85" *)
  wire _088_;
  (* src = "CanBtl.scala:141.43" *)
  wire _089_;
  (* src = "CanBtl.scala:141.40" *)
  wire _090_;
  (* src = "CanBtl.scala:141.95" *)
  wire [4:0] _091_;
  (* src = "CanBtl.scala:141.74" *)
  wire _092_;
  (* src = "CanBtl.scala:141.57" *)
  wire _093_;
  (* src = "CanBtl.scala:149.22" *)
  wire _094_;
  (* src = "CanBtl.scala:149.51" *)
  wire _095_;
  (* src = "CanBtl.scala:149.29" *)
  wire _096_;
  (* src = "CanBtl.scala:149.72" *)
  wire _097_;
  (* src = "CanBtl.scala:149.92" *)
  wire _098_;
  (* src = "CanBtl.scala:146.29" *)
  wire _099_;
  (* src = "CanBtl.scala:146.43" *)
  wire _100_;
  (* src = "CanBtl.scala:146.54" *)
  wire _101_;
  (* src = "CanBtl.scala:146.73" *)
  wire _102_;
  (* src = "CanBtl.scala:143.43" *)
  wire [6:0] _103_;
  (* src = "CanBtl.scala:143.43" *)
  wire [5:0] _104_;
  (* src = "CanBtl.scala:143.50" *)
  wire [6:0] _105_;
  (* src = "CanBtl.scala:197.36" *)
  wire [5:0] _106_;
  (* src = "CanBtl.scala:148.13" *)
  wire _107_;
  (* src = "CanBtl.scala:148.26" *)
  wire _108_;
  (* src = "CanBtl.scala:148.24" *)
  wire _109_;
  (* src = "CanBtl.scala:148.40" *)
  wire _110_;
  (* src = "CanBtl.scala:148.38" *)
  wire _111_;
  (* src = "CanBtl.scala:148.47" *)
  wire _112_;
  (* src = "CanBtl.scala:148.65" *)
  wire _113_;
  (* src = "CanBtl.scala:175.25" *)
  wire _114_;
  (* src = "Cat.scala:30.58" *)
  wire [1:0] _115_;
  (* src = "CanBtl.scala:214.34" *)
  wire _116_;
  (* src = "CanBtl.scala:214.50" *)
  wire _117_;
  (* src = "CanBtl.scala:214.37" *)
  wire _118_;
  (* src = "CanBtl.scala:214.68" *)
  wire _119_;
  (* src = "CanBtl.scala:214.72" *)
  wire _120_;
  (* src = "CanBtl.scala:214.59" *)
  wire _121_;
  (* src = "CanBtl.scala:151.50" *)
  wire [2:0] _122_;
  (* src = "CanBtl.scala:151.35" *)
  wire [3:0] _123_;
  (* src = "CanBtl.scala:151.35" *)
  wire [2:0] _124_;
  (* src = "CanBtl.scala:151.77" *)
  wire [4:0] _125_;
  (* src = "CanBtl.scala:151.77" *)
  wire [3:0] _126_;
  (* src = "CanBtl.scala:153.14" *)
  wire _127_;
  (* src = "CanBtl.scala:153.23" *)
  wire _128_;
  (* src = "CanBtl.scala:153.42" *)
  wire _129_;
  (* src = "CanBtl.scala:153.96" *)
  wire _130_;
  (* src = "CanBtl.scala:153.118" *)
  wire _131_;
  (* src = "CanBtl.scala:153.108" *)
  wire _132_;
  (* src = "CanBtl.scala:153.85" *)
  wire _133_;
  (* src = "CanBtl.scala:153.30" *)
  wire _134_;
  wire _135_;
  wire _136_;
  wire [1:0] _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire [6:0] _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  input clock;
  (* src = "CanBtl.scala:104.34" *)
  reg [6:0] clockCount;
  (* src = "CanBtl.scala:104.34|CanBtl.scala:104.34" *)
  wire [6:0] \clockCount$process$CanBtl_3 ;
  (* src = "CanBtl.scala:106.31" *)
  reg clockEn;
  (* src = "CanBtl.scala:106.31|CanBtl.scala:106.31" *)
  wire \clockEn$process$CanBtl_4 ;
  (* src = "CanBtl.scala:108.32" *)
  reg clockEnQ;
  (* src = "CanBtl.scala:108.32|CanBtl.scala:108.32|CanBtl.scala:108.32" *)
  wire \clockEnQ$process$CanBtl_5 ;
  (* src = "CanBtl.scala:116.29" *)
  reg [3:0] delay;
  (* src = "CanBtl.scala:116.29|CanBtl.scala:116.29" *)
  wire [3:0] \delay$process$CanBtl_9 ;
  (* src = "CanBtl.scala:138.32" *)
  wire goSeg1;
  (* src = "CanBtl.scala:141.32" *)
  wire goSeg2;
  (* src = "CanBtl.scala:149.89" *)
  wire goSync;
  (* src = "CanBtl.scala:112.39" *)
  reg hardSyncBlocked;
  (* src = "CanBtl.scala:112.39|CanBtl.scala:112.39" *)
  wire \hardSyncBlocked$process$CanBtl_7 ;
  input [5:0] io_baudRatePrescaler;
  input io_goErrorFrame;
  input io_goOverloadFrame;
  input io_goRxInter;
  input io_goTx;
  output io_hardSync;
  input io_nodeErrorPassive;
  input io_rx;
  input io_rxIdle;
  input io_rxInter;
  output io_samplePoint;
  output io_sampledBit;
  output io_sampledBitQ;
  input io_sendAck;
  input [1:0] io_syncJumpWidth;
  input [3:0] io_timeSegment1;
  input [2:0] io_timeSegment2;
  input io_transmitter;
  input io_transmitting;
  input io_tripleSampling;
  input io_tx;
  input io_txNext;
  output io_txPoint;
  (* src = "CanBtl.scala:132.35|CanBtl.scala:143.18" *)
  wire [7:0] prescalerLimit;
  (* src = "CanBtl.scala:114.37" *)
  reg [4:0] quantaCounter;
  (* src = "CanBtl.scala:114.37|CanBtl.scala:114.37" *)
  wire [4:0] \quantaCounter$process$CanBtl_8 ;
  input reset;
  (* src = "CanBtl.scala:148.63" *)
  wire resync;
  (* src = "CanBtl.scala:124.37" *)
  reg resyncLatched;
  (* src = "CanBtl.scala:124.37|CanBtl.scala:124.37" *)
  wire \resyncLatched$process$CanBtl_13 ;
  (* src = "CanBtl.scala:126.30" *)
  reg [1:0] sample;
  (* src = "CanBtl.scala:126.30|CanBtl.scala:126.30" *)
  wire [1:0] \sample$process$CanBtl_14 ;
  (* src = "CanBtl.scala:95.35" *)
  reg samplePoint;
  (* src = "CanBtl.scala:95.35|CanBtl.scala:95.35" *)
  wire \samplePoint$process$CanBtl ;
  (* src = "CanBtl.scala:99.34" *)
  reg sampledBit;
  (* src = "CanBtl.scala:99.34|CanBtl.scala:99.34" *)
  wire \sampledBit$process$CanBtl_1 ;
  (* src = "CanBtl.scala:101.35" *)
  reg sampledBitQ;
  (* src = "CanBtl.scala:101.35|CanBtl.scala:101.35" *)
  wire \sampledBitQ$process$CanBtl_2 ;
  (* src = "CanBtl.scala:120.28" *)
  reg seg1;
  (* src = "CanBtl.scala:120.28|CanBtl.scala:120.28" *)
  wire \seg1$process$CanBtl_11 ;
  (* src = "CanBtl.scala:122.28" *)
  reg seg2;
  (* src = "CanBtl.scala:122.28|CanBtl.scala:122.28" *)
  wire \seg2$process$CanBtl_12 ;
  (* src = "CanBtl.scala:118.28" *)
  reg sync;
  (* src = "CanBtl.scala:118.28|CanBtl.scala:118.28" *)
  wire \sync$process$CanBtl_10 ;
  (* src = "CanBtl.scala:110.35" *)
  reg syncBlocked;
  (* src = "CanBtl.scala:110.35|CanBtl.scala:110.35" *)
  wire \syncBlocked$process$CanBtl_6 ;
  (* src = "CanBtl.scala:151.57" *)
  wire syncWindow;
  (* src = "CanBtl.scala:128.31" *)
  reg txNextSp;
  (* src = "CanBtl.scala:128.31|CanBtl.scala:128.31" *)
  wire \txNextSp$process$CanBtl_15 ;
  (* src = "CanBtl.scala:97.31" *)
  reg txPoint;
  (* src = "CanBtl.scala:97.31|CanBtl.scala:97.31|CanBtl.scala:153.11" *)
  wire \txPoint$process$CanBtl_0 ;
  assign _125_ = { 1'h0, _025_ } + 5'h01;
  assign _091_ = { 1'h0, io_timeSegment1 } + { 1'h0, delay };
  assign _103_ = { 1'h0, io_baudRatePrescaler } + 7'h01;
  assign _079_ = { 1'h0, clockCount } + 8'h01;
  assign _106_ = { 1'h0, quantaCounter } + 6'h01;
  assign _109_ = _107_ & _108_;
  assign _111_ = _109_ & _110_;
  assign _112_ = _111_ & io_sampledBit;
  assign _100_ = _099_ & _110_;
  assign _101_ = _100_ & io_sampledBit;
  assign _094_ = clockEnQ & seg2;
  assign _096_ = _094_ & _095_;
  assign _097_ = _096_ & _089_;
  assign goSync = _097_ & _098_;
  assign _128_ = _127_ & seg2;
  assign _129_ = clockEn & _095_;
  assign _132_ = _130_ & _131_;
  assign _134_ = _128_ & _133_;
  assign resync = _112_ & _113_;
  assign _077_ = _084_ & _076_;
  assign _049_ = resync & seg1;
  assign _051_ = io_tx & _110_;
  assign _053_ = io_transmitting & _052_;
  assign _055_ = _049_ & _054_;
  assign _057_ = clockEnQ & _089_;
  assign _058_ = seg1 & _092_;
  assign _117_ = _114_ & io_rx;
  assign _120_ = _119_ & io_rx;
  assign _010_ = _057_ & _007_;
  assign _084_ = resync & seg2;
  assign _060_ = io_goErrorFrame & _059_;
  assign _064_ = io_goErrorFrame & io_nodeErrorPassive;
  assign _065_ = io_hardSync & clockEnQ;
  assign _066_ = io_transmitting & io_transmitter;
  assign _068_ = _067_ & io_txPoint;
  assign _070_ = _068_ & _069_;
  assign _072_ = _099_ & samplePoint;
  assign _073_ = _072_ & io_sampledBit;
  assign io_hardSync = _101_ & _102_;
  assign _085_ = _084_ & syncWindow;
  assign _087_ = resyncLatched & syncWindow;
  assign goSeg1 = clockEnQ & _088_;
  assign _090_ = seg1 & _089_;
  assign _093_ = _090_ & _092_;
  assign goSeg2 = clockEnQ & _093_;
  assign _092_ = quantaCounter == _091_;
  assign _095_ = _122_ == io_timeSegment2;
  assign _075_ = _027_ == _047_;
  assign _056_ = _027_ >= _047_;
  assign _081_ = quantaCounter > _028_;
  assign syncWindow = _026_ < _126_;
  assign _000_ = _056_ ? (* src = "CanBtl.scala:155.46|CanBtl.scala:156.16|CanBtl.scala:158.16" *) 7'h00 : _080_;
  assign _011_ = goSeg1 ? (* src = "CanBtl.scala:169.22|CanBtl.scala:170.19|CanBtl.scala:124.37" *) 1'h0 : resyncLatched;
  assign _031_ = clockEnQ ? (* src = "CanBtl.scala:173.18|CanBtl.scala:174.10|CanBtl.scala:118.28" *) goSync : sync;
  assign _005_ = io_tripleSampling ? (* src = "CanBtl.scala:213.31|CanBtl.scala:214.20|CanBtl.scala:216.20" *) _121_ : io_rx;
  assign _006_ = _058_ ? (* src = "CanBtl.scala:212.65|CanBtl.scala:99.34" *) _005_ : sampledBit;
  assign _008_ = _058_ ? (* src = "CanBtl.scala:212.65|CanBtl.scala:219.19|CanBtl.scala:101.35" *) sampledBit : sampledBitQ;
  assign _009_ = _057_ ? (* src = "CanBtl.scala:211.38|CanBtl.scala:99.34" *) _006_ : sampledBit;
  assign _012_ = _057_ ? (* src = "CanBtl.scala:211.38|CanBtl.scala:101.35" *) _008_ : sampledBitQ;
  assign _013_ = io_goErrorFrame ? (* src = "CanBtl.scala:207.25|CanBtl.scala:208.17" *) sampledBit : _012_;
  assign _014_ = io_goErrorFrame ? (* src = "CanBtl.scala:207.25|CanBtl.scala:209.17" *) 1'h0 : _010_;
  assign _015_ = io_goErrorFrame ? (* src = "CanBtl.scala:207.25|CanBtl.scala:99.34" *) sampledBit : _009_;
  assign _016_ = samplePoint ? (* src = "CanBtl.scala:231.26|CanBtl.scala:232.14|CanBtl.scala:128.31" *) io_txNext : txNextSp;
  assign _018_ = _063_ ? (* src = "CanBtl.scala:225.94|CanBtl.scala:226.14" *) 1'h0 : _017_;
  assign _032_ = clockEnQ ? (* src = "CanBtl.scala:173.18|CanBtl.scala:175.12|CanBtl.scala:126.30" *) _115_ : sample;
  assign _019_ = goSeg2 ? (* src = "CanBtl.scala:238.24|CanBtl.scala:239.19|CanBtl.scala:110.35" *) 1'h0 : syncBlocked;
  assign _021_ = clockEnQ ? (* src = "CanBtl.scala:235.18|CanBtl.scala:110.35" *) _020_ : syncBlocked;
  assign _023_ = _074_ ? (* src = "CanBtl.scala:246.84|CanBtl.scala:247.21|CanBtl.scala:112.39" *) 1'h0 : hardSyncBlocked;
  assign _029_ = reset ? (* src = "CanBtl.scala:114.37|CanBtl.scala:114.37" *) 6'h00 : _002_;
  assign _030_ = reset ? (* src = "CanBtl.scala:116.29|CanBtl.scala:116.29" *) 6'h00 : _004_;
  assign _033_ = goSeg2 ? (* src = "CanBtl.scala:181.22|CanBtl.scala:183.10|CanBtl.scala:120.28" *) 1'h0 : seg1;
  assign _035_ = _078_ ? (* src = "CanBtl.scala:188.31|CanBtl.scala:189.10|CanBtl.scala:122.28" *) 1'h0 : seg2;
  assign _001_ = clockEnQ ? (* src = "CanBtl.scala:195.24|CanBtl.scala:197.19|CanBtl.scala:114.37" *) _106_ : { 1'h0, quantaCounter };
  assign _002_ = _048_ ? (* src = "CanBtl.scala:192.34|CanBtl.scala:194.19" *) 6'h00 : _001_;
  assign _082_ = _081_ ? (* src = "CanBtl.scala:201.17" *) { 2'h0, _126_ } : _106_;
  assign _003_ = _078_ ? (* src = "CanBtl.scala:203.30|CanBtl.scala:204.11|CanBtl.scala:116.29" *) 4'h0 : delay;
  assign _004_ = _055_ ? (* src = "CanBtl.scala:200.94|CanBtl.scala:201.11" *) _082_ : { 2'h0, _003_ };
  assign _107_ = ~ io_rxIdle;
  assign _108_ = ~ io_rxInter;
  assign _110_ = ~ io_rx;
  assign _069_ = ~ io_txNext;
  assign _113_ = ~ syncBlocked;
  assign _089_ = ~ io_hardSync;
  assign _102_ = ~ hardSyncBlocked;
  assign _098_ = ~ resync;
  assign _127_ = ~ txPoint;
  assign _076_ = ~ syncWindow;
  assign _050_ = ~ io_transmitting;
  assign _059_ = ~ io_nodeErrorPassive;
  assign _037_ = reset | _015_;
  assign _038_ = reset | _013_;
  assign _039_ = reset | _021_;
  assign _022_ = _077_ | _011_;
  assign _034_ = goSeg1 | _033_;
  assign _078_ = goSync | goSeg1;
  assign _036_ = goSeg2 | _035_;
  assign _048_ = _078_ | goSeg2;
  assign _052_ = txNextSp | _051_;
  assign _054_ = _050_ | _053_;
  assign _118_ = _116_ | _117_;
  assign _121_ = _118_ | _120_;
  assign _007_ = _058_ | samplePoint;
  assign _042_ = reset | _034_;
  assign _061_ = io_goOverloadFrame | _060_;
  assign _062_ = _061_ | io_goTx;
  assign _063_ = _062_ | io_sendAck;
  assign _017_ = _064_ | _016_;
  assign _020_ = resync | _019_;
  assign _067_ = _066_ | io_goTx;
  assign _071_ = _065_ | _070_;
  assign _074_ = io_goRxInter | _073_;
  assign _024_ = _071_ | _023_;
  assign _083_ = sync | io_hardSync;
  assign _086_ = _083_ | _085_;
  assign _088_ = _086_ | _087_;
  assign _099_ = io_rxIdle | io_rxInter;
  assign _130_ = clockEn | clockEnQ;
  assign _131_ = resync | io_hardSync;
  assign _133_ = _129_ | _132_;
  always @(posedge clock)
    txNextSp <= _135_;
  always @(posedge clock)
    sample <= _137_;
  always @(posedge clock)
    resyncLatched <= _139_;
  always @(posedge clock)
    seg2 <= _141_;
  always @(posedge clock)
    seg1 <= _042_;
  always @(posedge clock)
    sync <= _143_;
  always @(posedge clock)
    delay <= _030_[3:0];
  always @(posedge clock)
    quantaCounter <= _029_[4:0];
  always @(posedge clock)
    hardSyncBlocked <= _145_;
  always @(posedge clock)
    syncBlocked <= _039_;
  always @(posedge clock)
    clockEnQ <= _147_;
  always @(posedge clock)
    clockEn <= _149_;
  always @(posedge clock)
    clockCount <= _151_;
  always @(posedge clock)
    sampledBitQ <= _038_;
  always @(posedge clock)
    sampledBit <= _037_;
  always @(posedge clock)
    txPoint <= _153_;
  always @(posedge clock)
    samplePoint <= _155_;
  assign _135_ = _136_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:128.31" *) 1'h0 : _018_;
  assign _137_ = _138_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:126.30" *) 2'h3 : _032_;
  assign _139_ = _140_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:124.37" *) 1'h0 : _022_;
  assign _141_ = _142_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:122.28" *) 1'h0 : _036_;
  assign _143_ = _144_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:118.28" *) 1'h0 : _031_;
  assign _145_ = _146_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:112.39" *) 1'h0 : _024_;
  assign _147_ = _148_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:108.32" *) 1'h0 : clockEn;
  assign _149_ = _150_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:106.31" *) 1'h0 : _075_;
  assign _151_ = _152_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:104.34" *) 7'h00 : _000_;
  assign _153_ = _154_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:97.31" *) 1'h0 : _134_;
  assign _155_ = _156_ ? (* full_case = 32'd1 *) (* src = "CanBtl.scala:95.35" *) 1'h0 : _014_;
  assign _116_ = & sample;
  assign _123_ = { 1'h0, io_timeSegment2 } - { 1'h0, _122_ };
  assign _046_ = { 1'h0, prescalerLimit } - 9'h001;
  assign _122_ = quantaCounter[2:0];
  assign _124_ = _123_[2:0];
  assign _025_ = { 2'h0, io_syncJumpWidth };
  assign _126_ = _125_[3:0];
  assign _026_ = { 1'h0, _124_ };
  assign _104_ = _103_[5:0];
  assign _105_ = { _104_, 1'h0 };
  assign prescalerLimit = { 1'h0, _105_ };
  assign _047_ = _046_[7:0];
  assign _027_ = { 1'h0, clockCount };
  assign _080_ = _079_[6:0];
  assign _114_ = sample[0];
  assign _115_ = { _114_, io_rx };
  assign _028_ = { 3'h0, io_syncJumpWidth };
  assign _119_ = sample[1];
  assign io_samplePoint = samplePoint;
  assign io_sampledBit = sampledBit;
  assign io_sampledBitQ = sampledBitQ;
  assign io_txPoint = txPoint;
  assign \seg1$process$CanBtl_11  = _042_;
  assign \delay$process$CanBtl_9  = _030_[3:0];
  assign \quantaCounter$process$CanBtl_8  = _029_[4:0];
  assign \syncBlocked$process$CanBtl_6  = _039_;
  assign \sampledBitQ$process$CanBtl_2  = _038_;
  assign \sampledBit$process$CanBtl_1  = _037_;
  assign _136_ = reset;
  assign \txNextSp$process$CanBtl_15  = _135_;
  assign _138_ = reset;
  assign \sample$process$CanBtl_14  = _137_;
  assign _140_ = reset;
  assign \resyncLatched$process$CanBtl_13  = _139_;
  assign _142_ = reset;
  assign \seg2$process$CanBtl_12  = _141_;
  assign _144_ = reset;
  assign \sync$process$CanBtl_10  = _143_;
  assign _146_ = reset;
  assign \hardSyncBlocked$process$CanBtl_7  = _145_;
  assign _148_ = reset;
  assign \clockEnQ$process$CanBtl_5  = _147_;
  assign _150_ = reset;
  assign \clockEn$process$CanBtl_4  = _149_;
  assign _152_ = reset;
  assign \clockCount$process$CanBtl_3  = _151_;
  assign _154_ = reset;
  assign \txPoint$process$CanBtl_0  = _153_;
  assign _156_ = reset;
  assign \samplePoint$process$CanBtl  = _155_;
endmodule

(* cells_not_processed =  1  *)
module CanCrc(clock, reset, io_data, io_enable, io_crc);
  (* src = "CanCrc.scala:19.19|CanCrc.scala:20.11|CanCrc.scala:22.11" *)
  wire [14:0] _00_;
  (* src = "CanCrc.scala:18.19|CanCrc.scala:13.27" *)
  wire [14:0] _01_;
  (* src = "CanCrc.scala:14.40" *)
  wire _02_;
  (* src = "CanCrc.scala:15.33" *)
  wire [13:0] _03_;
  (* src = "CanCrc.scala:20.21" *)
  wire [14:0] _04_;
  wire [14:0] _05_;
  wire _06_;
  input clock;
  (* src = "CanCrc.scala:13.27" *)
  reg [14:0] crc;
  (* src = "CanCrc.scala:13.27|CanCrc.scala:13.27" *)
  wire [14:0] \crc$process$CanCrc ;
  (* src = "CanCrc.scala:14.32" *)
  wire crcNext;
  (* src = "Cat.scala:30.58" *)
  wire [14:0] crcTmp;
  output [14:0] io_crc;
  input io_data;
  input io_enable;
  input reset;
  assign _00_ = crcNext ? (* src = "CanCrc.scala:19.19|CanCrc.scala:20.11|CanCrc.scala:22.11" *) _04_ : crcTmp;
  assign _01_ = io_enable ? (* src = "CanCrc.scala:18.19|CanCrc.scala:13.27" *) _00_ : crc;
  always @(posedge clock)
    crc <= _05_;
  assign _05_ = _06_ ? (* full_case = 32'd1 *) (* src = "CanCrc.scala:13.27" *) 15'h0000 : _01_;
  assign crcNext = io_data ^ _02_;
  assign _04_ = crcTmp ^ 15'h4599;
  assign _02_ = io_crc[14];
  assign _03_ = io_crc[13:0];
  assign crcTmp = { _03_, 1'h0 };
  assign io_crc = crc;
  assign _06_ = reset;
  assign \crc$process$CanCrc  = _05_;
endmodule

(* cells_not_processed =  1  *)
module CanFifo(clock, reset, io_wr, io_dataIn, io_addr, io_dataOut, io_resetMode, io_releaseBuffer, io_extendedMode, io_overrun, io_infoEmpty, io_infoCnt);
  (* src = "CanFifo.scala:63.35|CanFifo.scala:64.12|CanFifo.scala:47.30" *)
  wire [3:0] _000_;
  (* src = "CanFifo.scala:61.40|CanFifo.scala:62.12" *)
  wire [3:0] _001_;
  (* src = "CanFifo.scala:87.40|CanFifo.scala:88.18" *)
  wire _002_;
  (* src = "CanFifo.scala:99.65|CanFifo.scala:100.15|CanFifo.scala:48.31" *)
  wire [7:0] _003_;
  (* src = "CanFifo.scala:97.54|CanFifo.scala:98.13" *)
  wire [7:0] _004_;
  (* src = "CanFifo.scala:95.53|CanFifo.scala:96.13" *)
  wire [7:0] _005_;
  (* src = "CanFifo.scala:93.22|CanFifo.scala:94.13" *)
  wire [7:0] _006_;
  (* src = "CanFifo.scala:108.45|CanFifo.scala:109.15|CanFifo.scala:23.31" *)
  wire [7:0] _007_;
  (* src = "CanFifo.scala:106.44|CanFifo.scala:107.15" *)
  wire [7:0] _008_;
  (* src = "CanFifo.scala:105.50|CanFifo.scala:23.31" *)
  wire [7:0] _009_;
  (* src = "CanFifo.scala:103.22|CanFifo.scala:104.13" *)
  wire [7:0] _010_;
  (* src = "CanFifo.scala:113.30|CanFifo.scala:114.24|CanFifo.scala:51.42" *)
  wire _011_;
  (* src = "CanFifo.scala:69.28|CanFifo.scala:70.19|CanFifo.scala:44.37" *)
  wire [5:0] _012_;
  (* src = "CanFifo.scala:67.60|CanFifo.scala:68.19" *)
  wire [5:0] _013_;
  (* src = "CanFifo.scala:78.28" *)
  wire [5:0] _014_;
  (* src = "CanFifo.scala:23.31|CanFifo.scala:23.31" *)
  wire [7:0] _015_;
  (* src = "CanFifo.scala:45.37|CanFifo.scala:45.37" *)
  wire [6:0] _016_;
  (* src = "CanFifo.scala:48.31|CanFifo.scala:48.31" *)
  wire [7:0] _017_;
  (* src = "CanFifo.scala:73.38|CanFifo.scala:74.19|CanFifo.scala:45.37" *)
  wire [6:0] _018_;
  (* src = "CanFifo.scala:77.39|CanFifo.scala:78.15|CanFifo.scala:41.33" *)
  wire [5:0] _019_;
  (* src = "CanFifo.scala:83.33|CanFifo.scala:84.15|CanFifo.scala:42.33" *)
  wire [5:0] _020_;
  (* src = "CanFifo.scala:81.22|CanFifo.scala:82.15" *)
  wire [5:0] _021_;
  (* src = "CanFifo.scala:89.32|CanFifo.scala:90.18|CanFifo.scala:50.36" *)
  wire _022_;
  wire [5:0] _023_;
  wire [3:0] _024_;
  wire _025_;
  wire _026_;
  wire [7:0] _027_;
  wire [7:0] _028_;
  wire [7:0] _029_;
  wire [7:0] _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire [6:0] _034_;
  wire [5:0] _035_;
  wire [6:0] _036_;
  wire _037_;
  wire [6:0] _038_;
  (* src = "CanFifo.scala:61.21" *)
  wire _039_;
  (* src = "CanFifo.scala:63.23" *)
  wire _040_;
  (* src = "CanFifo.scala:89.20" *)
  wire _041_;
  (* src = "CanFifo.scala:95.22" *)
  wire _042_;
  (* src = "CanFifo.scala:95.20" *)
  wire _043_;
  (* src = "CanFifo.scala:95.40" *)
  wire _044_;
  (* src = "CanFifo.scala:97.21" *)
  wire _045_;
  (* src = "CanFifo.scala:63.20" *)
  wire _046_;
  (* src = "CanFifo.scala:97.40" *)
  wire _047_;
  (* src = "CanFifo.scala:99.20" *)
  wire _048_;
  (* src = "CanFifo.scala:99.39" *)
  wire _049_;
  (* src = "CanFifo.scala:99.51" *)
  wire _050_;
  (* src = "CanFifo.scala:105.30" *)
  wire _051_;
  (* src = "CanFifo.scala:106.29" *)
  wire _052_;
  (* src = "CanFifo.scala:106.27" *)
  wire _053_;
  (* src = "CanFifo.scala:67.27" *)
  wire _054_;
  (* src = "CanFifo.scala:113.26" *)
  wire _055_;
  (* src = "CanFifo.scala:67.24" *)
  wire _056_;
  (* src = "CanFifo.scala:128.51" *)
  wire _057_;
  (* src = "CanFifo.scala:128.76" *)
  wire _058_;
  (* src = "CanFifo.scala:67.38" *)
  wire _059_;
  (* src = "CanFifo.scala:73.25" *)
  wire _060_;
  (* src = "CanFifo.scala:77.27" *)
  wire _061_;
  (* src = "CanFifo.scala:77.25" *)
  wire _062_;
  (* src = "CanFifo.scala:96.24" *)
  wire [7:0] _063_;
  (* src = "Cat.scala:30.58" *)
  wire [6:0] _064_;
  (* src = "CanFifo.scala:98.24" *)
  wire [7:0] _065_;
  (* src = "CanFifo.scala:98.24" *)
  wire [6:0] _066_;
  (* src = "CanFifo.scala:100.53" *)
  wire [7:0] _067_;
  (* src = "CanFifo.scala:107.27" *)
  wire [7:0] _068_;
  (* src = "CanFifo.scala:109.27" *)
  wire [7:0] _069_;
  (* src = "CanFifo.scala:64.22" *)
  wire [4:0] _070_;
  (* src = "CanFifo.scala:64.22" *)
  wire [3:0] _071_;
  (* src = "CanFifo.scala:74.36" *)
  wire [6:0] _072_;
  (* src = "CanFifo.scala:78.28" *)
  wire [6:0] _073_;
  (* src = "CanFifo.scala:78.28" *)
  wire [5:0] _074_;
  (* src = "CanFifo.scala:59.45" *)
  wire [5:0] _075_;
  (* src = "CanFifo.scala:59.40" *)
  wire [6:0] _076_;
  (* src = "CanFifo.scala:59.40" *)
  wire [5:0] _077_;
  (* src = "CanFifo.scala:59.29" *)
  wire [6:0] _078_;
  (* src = "CanFifo.scala:68.36" *)
  wire [6:0] _079_;
  (* src = "CanFifo.scala:68.36" *)
  wire [5:0] _080_;
  (* src = "CanFifo.scala:84.28" *)
  wire [6:0] _081_;
  (* src = "CanFifo.scala:84.28" *)
  wire [5:0] _082_;
  (* src = "CanFifo.scala:46.31" *)
  wire _083_;
  (* src = "CanFifo.scala:53.32" *)
  wire _084_;
  wire [7:0] _085_;
  wire [3:0] _086_;
  wire _087_;
  wire _088_;
  wire [3:0] _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire [5:0] _093_;
  wire _094_;
  wire [5:0] _095_;
  wire _096_;
  wire [5:0] _097_;
  wire _098_;
  input clock;
  (* src = "CanFifo.scala:48.31" *)
  reg [6:0] fifoCnt;
  (* src = "CanFifo.scala:48.31|CanFifo.scala:48.31" *)
  wire [6:0] \fifoCnt$process$CanFifo_6 ;
  (* src = "CanFifo.scala:54.34" *)
  wire fifoEmpty;
  (* src = "CanFifo.scala:55.33" *)
  wire fifoFull;
  wire [7:0] fifo_io_dataOut_MPORT_data;
  (* src = "CanFifo.scala:23.31" *)
  reg [6:0] infoCnt;
  (* src = "CanFifo.scala:23.31|CanFifo.scala:23.31" *)
  wire [6:0] \infoCnt$process$CanFifo ;
  (* src = "CanFifo.scala:56.33" *)
  wire infoFull;
  (* src = "CanFifo.scala:51.42" *)
  reg initializeMemories;
  (* src = "CanFifo.scala:51.42|CanFifo.scala:51.42" *)
  wire \initializeMemories$process$CanFifo_8 ;
  input [5:0] io_addr;
  input [7:0] io_dataIn;
  output [7:0] io_dataOut;
  input io_extendedMode;
  output [6:0] io_infoCnt;
  output io_infoEmpty;
  output io_overrun;
  input io_releaseBuffer;
  input io_resetMode;
  input io_wr;
  (* src = "CanFifo.scala:50.36" *)
  reg latchOverrun;
  (* src = "CanFifo.scala:50.36|CanFifo.scala:50.36" *)
  wire \latchOverrun$process$CanFifo_7 ;
  (* src = "CanFifo.scala:47.30" *)
  reg [3:0] lenCnt;
  (* src = "CanFifo.scala:47.30|CanFifo.scala:47.30" *)
  wire [3:0] \lenCnt$process$CanFifo_5 ;
  wire [3:0] lengthFifo_lengthInfo_MPORT_data;
  (* src = "CanFifo.scala:52.31|CanFifo.scala:58.14" *)
  wire [3:0] lengthInfo;
  wire overrunInfo_io_overrun_MPORT_data;
  (* src = "CanFifo.scala:45.37" *)
  reg [5:0] rdInfoPointer;
  (* src = "CanFifo.scala:45.37|CanFifo.scala:45.37" *)
  wire [5:0] \rdInfoPointer$process$CanFifo_3 ;
  (* src = "CanFifo.scala:41.33" *)
  reg [5:0] rdPointer;
  (* src = "CanFifo.scala:41.33|CanFifo.scala:41.33" *)
  wire [5:0] \rdPointer$process$CanFifo_0 ;
  input reset;
  (* src = "CanFifo.scala:44.37" *)
  reg [5:0] wrInfoPointer;
  (* src = "CanFifo.scala:44.37|CanFifo.scala:44.37" *)
  wire [5:0] \wrInfoPointer$process$CanFifo_2 ;
  (* src = "CanFifo.scala:42.33" *)
  reg [5:0] wrPointer;
  (* src = "CanFifo.scala:42.33|CanFifo.scala:42.33" *)
  wire [5:0] \wrPointer$process$CanFifo_1 ;
  (* src = "CanFifo.scala:46.27" *)
  reg wrQ;
  (* src = "CanFifo.scala:46.27|CanFifo.scala:46.27|CanFifo.scala:46.27" *)
  wire \wrQ$process$CanFifo_4 ;
  (* src = "CanFifo.scala:53.39" *)
  wire writeLengthInfo;
  reg [7:0] fifo [63:0];
  initial begin
    fifo[0] = 8'h00;
    fifo[1] = 8'h00;
    fifo[2] = 8'h00;
    fifo[3] = 8'h00;
    fifo[4] = 8'h00;
    fifo[5] = 8'h00;
    fifo[6] = 8'h00;
    fifo[7] = 8'h00;
    fifo[8] = 8'h00;
    fifo[9] = 8'h00;
    fifo[10] = 8'h00;
    fifo[11] = 8'h00;
    fifo[12] = 8'h00;
    fifo[13] = 8'h00;
    fifo[14] = 8'h00;
    fifo[15] = 8'h00;
    fifo[16] = 8'h00;
    fifo[17] = 8'h00;
    fifo[18] = 8'h00;
    fifo[19] = 8'h00;
    fifo[20] = 8'h00;
    fifo[21] = 8'h00;
    fifo[22] = 8'h00;
    fifo[23] = 8'h00;
    fifo[24] = 8'h00;
    fifo[25] = 8'h00;
    fifo[26] = 8'h00;
    fifo[27] = 8'h00;
    fifo[28] = 8'h00;
    fifo[29] = 8'h00;
    fifo[30] = 8'h00;
    fifo[31] = 8'h00;
    fifo[32] = 8'h00;
    fifo[33] = 8'h00;
    fifo[34] = 8'h00;
    fifo[35] = 8'h00;
    fifo[36] = 8'h00;
    fifo[37] = 8'h00;
    fifo[38] = 8'h00;
    fifo[39] = 8'h00;
    fifo[40] = 8'h00;
    fifo[41] = 8'h00;
    fifo[42] = 8'h00;
    fifo[43] = 8'h00;
    fifo[44] = 8'h00;
    fifo[45] = 8'h00;
    fifo[46] = 8'h00;
    fifo[47] = 8'h00;
    fifo[48] = 8'h00;
    fifo[49] = 8'h00;
    fifo[50] = 8'h00;
    fifo[51] = 8'h00;
    fifo[52] = 8'h00;
    fifo[53] = 8'h00;
    fifo[54] = 8'h00;
    fifo[55] = 8'h00;
    fifo[56] = 8'h00;
    fifo[57] = 8'h00;
    fifo[58] = 8'h00;
    fifo[59] = 8'h00;
    fifo[60] = 8'h00;
    fifo[61] = 8'h00;
    fifo[62] = 8'h00;
    fifo[63] = 8'h00;
  end
  always @(posedge clock) begin
    if (_085_[0])
      fifo[wrPointer][0:0] <= io_dataIn[0];
    if (_085_[1])
      fifo[wrPointer][1:1] <= io_dataIn[1];
    if (_085_[2])
      fifo[wrPointer][2:2] <= io_dataIn[2];
    if (_085_[3])
      fifo[wrPointer][3:3] <= io_dataIn[3];
    if (_085_[4])
      fifo[wrPointer][4:4] <= io_dataIn[4];
    if (_085_[5])
      fifo[wrPointer][5:5] <= io_dataIn[5];
    if (_085_[6])
      fifo[wrPointer][6:6] <= io_dataIn[6];
    if (_085_[7])
      fifo[wrPointer][7:7] <= io_dataIn[7];
  end
  reg [7:0] _388_;
  always @(posedge clock) begin
    _388_ <= fifo[_078_[5:0]];
  end
  assign fifo_io_dataOut_MPORT_data = _388_;
  reg [3:0] lengthFifo [63:0];
  initial begin
    lengthFifo[0] = 4'h0;
    lengthFifo[1] = 4'h0;
    lengthFifo[2] = 4'h0;
    lengthFifo[3] = 4'h0;
    lengthFifo[4] = 4'h0;
    lengthFifo[5] = 4'h0;
    lengthFifo[6] = 4'h0;
    lengthFifo[7] = 4'h0;
    lengthFifo[8] = 4'h0;
    lengthFifo[9] = 4'h0;
    lengthFifo[10] = 4'h0;
    lengthFifo[11] = 4'h0;
    lengthFifo[12] = 4'h0;
    lengthFifo[13] = 4'h0;
    lengthFifo[14] = 4'h0;
    lengthFifo[15] = 4'h0;
    lengthFifo[16] = 4'h0;
    lengthFifo[17] = 4'h0;
    lengthFifo[18] = 4'h0;
    lengthFifo[19] = 4'h0;
    lengthFifo[20] = 4'h0;
    lengthFifo[21] = 4'h0;
    lengthFifo[22] = 4'h0;
    lengthFifo[23] = 4'h0;
    lengthFifo[24] = 4'h0;
    lengthFifo[25] = 4'h0;
    lengthFifo[26] = 4'h0;
    lengthFifo[27] = 4'h0;
    lengthFifo[28] = 4'h0;
    lengthFifo[29] = 4'h0;
    lengthFifo[30] = 4'h0;
    lengthFifo[31] = 4'h0;
    lengthFifo[32] = 4'h0;
    lengthFifo[33] = 4'h0;
    lengthFifo[34] = 4'h0;
    lengthFifo[35] = 4'h0;
    lengthFifo[36] = 4'h0;
    lengthFifo[37] = 4'h0;
    lengthFifo[38] = 4'h0;
    lengthFifo[39] = 4'h0;
    lengthFifo[40] = 4'h0;
    lengthFifo[41] = 4'h0;
    lengthFifo[42] = 4'h0;
    lengthFifo[43] = 4'h0;
    lengthFifo[44] = 4'h0;
    lengthFifo[45] = 4'h0;
    lengthFifo[46] = 4'h0;
    lengthFifo[47] = 4'h0;
    lengthFifo[48] = 4'h0;
    lengthFifo[49] = 4'h0;
    lengthFifo[50] = 4'h0;
    lengthFifo[51] = 4'h0;
    lengthFifo[52] = 4'h0;
    lengthFifo[53] = 4'h0;
    lengthFifo[54] = 4'h0;
    lengthFifo[55] = 4'h0;
    lengthFifo[56] = 4'h0;
    lengthFifo[57] = 4'h0;
    lengthFifo[58] = 4'h0;
    lengthFifo[59] = 4'h0;
    lengthFifo[60] = 4'h0;
    lengthFifo[61] = 4'h0;
    lengthFifo[62] = 4'h0;
    lengthFifo[63] = 4'h0;
  end
  always @(posedge clock) begin
    if (_086_[0])
      lengthFifo[wrInfoPointer][0:0] <= _024_[0];
    if (_086_[1])
      lengthFifo[wrInfoPointer][1:1] <= _024_[1];
    if (_086_[2])
      lengthFifo[wrInfoPointer][2:2] <= _024_[2];
    if (_086_[3])
      lengthFifo[wrInfoPointer][3:3] <= _024_[3];
  end
  reg [3:0] _389_;
  always @(posedge clock) begin
    if (1'h0) begin
      _389_ <= lengthFifo[rdInfoPointer];
    end
  end
  assign lengthFifo_lengthInfo_MPORT_data = _389_;
  reg [0:0] overrunInfo [63:0];
  initial begin
    overrunInfo[0] = 1'h0;
    overrunInfo[1] = 1'h0;
    overrunInfo[2] = 1'h0;
    overrunInfo[3] = 1'h0;
    overrunInfo[4] = 1'h0;
    overrunInfo[5] = 1'h0;
    overrunInfo[6] = 1'h0;
    overrunInfo[7] = 1'h0;
    overrunInfo[8] = 1'h0;
    overrunInfo[9] = 1'h0;
    overrunInfo[10] = 1'h0;
    overrunInfo[11] = 1'h0;
    overrunInfo[12] = 1'h0;
    overrunInfo[13] = 1'h0;
    overrunInfo[14] = 1'h0;
    overrunInfo[15] = 1'h0;
    overrunInfo[16] = 1'h0;
    overrunInfo[17] = 1'h0;
    overrunInfo[18] = 1'h0;
    overrunInfo[19] = 1'h0;
    overrunInfo[20] = 1'h0;
    overrunInfo[21] = 1'h0;
    overrunInfo[22] = 1'h0;
    overrunInfo[23] = 1'h0;
    overrunInfo[24] = 1'h0;
    overrunInfo[25] = 1'h0;
    overrunInfo[26] = 1'h0;
    overrunInfo[27] = 1'h0;
    overrunInfo[28] = 1'h0;
    overrunInfo[29] = 1'h0;
    overrunInfo[30] = 1'h0;
    overrunInfo[31] = 1'h0;
    overrunInfo[32] = 1'h0;
    overrunInfo[33] = 1'h0;
    overrunInfo[34] = 1'h0;
    overrunInfo[35] = 1'h0;
    overrunInfo[36] = 1'h0;
    overrunInfo[37] = 1'h0;
    overrunInfo[38] = 1'h0;
    overrunInfo[39] = 1'h0;
    overrunInfo[40] = 1'h0;
    overrunInfo[41] = 1'h0;
    overrunInfo[42] = 1'h0;
    overrunInfo[43] = 1'h0;
    overrunInfo[44] = 1'h0;
    overrunInfo[45] = 1'h0;
    overrunInfo[46] = 1'h0;
    overrunInfo[47] = 1'h0;
    overrunInfo[48] = 1'h0;
    overrunInfo[49] = 1'h0;
    overrunInfo[50] = 1'h0;
    overrunInfo[51] = 1'h0;
    overrunInfo[52] = 1'h0;
    overrunInfo[53] = 1'h0;
    overrunInfo[54] = 1'h0;
    overrunInfo[55] = 1'h0;
    overrunInfo[56] = 1'h0;
    overrunInfo[57] = 1'h0;
    overrunInfo[58] = 1'h0;
    overrunInfo[59] = 1'h0;
    overrunInfo[60] = 1'h0;
    overrunInfo[61] = 1'h0;
    overrunInfo[62] = 1'h0;
    overrunInfo[63] = 1'h0;
  end
  always @(posedge clock) begin
    if (_032_)
      overrunInfo[wrInfoPointer] <= _033_;
  end
  reg [0:0] _390_;
  always @(posedge clock) begin
    if (_031_) begin
      _390_ <= overrunInfo[rdInfoPointer];
    end
  end
  assign overrunInfo_io_overrun_MPORT_data = _390_;
  assign _078_ = { 1'h0, rdPointer } + { 1'h0, _077_ };
  assign _070_ = { 1'h0, lenCnt } + 5'h01;
  assign _079_ = { 1'h0, wrInfoPointer } + 7'h01;
  assign _072_ = { 1'h0, rdInfoPointer } + 7'h01;
  assign _073_ = { 1'h0, rdPointer } + { 1'h0, _014_ };
  assign _081_ = { 1'h0, wrPointer } + 7'h01;
  assign _063_ = { 1'h0, fifoCnt } + 8'h01;
  assign _067_ = { 1'h0, _066_ } + 8'h01;
  assign _069_ = { 1'h0, infoCnt } + 8'h01;
  assign _025_ = io_wr & _040_;
  assign _085_ = $signed(_025_) & (* src = "CanFifo.scala:37.45" *) $signed(1'h1);
  assign _086_ = $signed(_026_) & (* src = "CanFifo.scala:38.51" *) $signed(1'h1);
  assign _043_ = io_wr & _042_;
  assign _044_ = _043_ & _040_;
  assign _045_ = _084_ & io_releaseBuffer;
  assign _047_ = _045_ & _061_;
  assign _048_ = io_wr & io_releaseBuffer;
  assign _049_ = _048_ & _040_;
  assign _050_ = _049_ & _061_;
  assign _053_ = io_releaseBuffer & _052_;
  assign _031_ = io_releaseBuffer & _054_;
  assign _033_ = _057_ & _058_;
  assign writeLengthInfo = _084_ & wrQ;
  assign _046_ = io_wr & _040_;
  assign _056_ = writeLengthInfo & _054_;
  assign _060_ = io_releaseBuffer & _054_;
  assign _062_ = io_releaseBuffer & _061_;
  assign _041_ = io_wr & fifoFull;
  assign fifoEmpty = ! fifoCnt;
  assign fifoFull = fifoCnt == 7'h40;
  assign infoFull = infoCnt == 7'h40;
  assign io_infoEmpty = ! infoCnt;
  assign _024_ = initializeMemories ? (* src = "CanFifo.scala:124.37" *) 4'h0 : lenCnt;
  assign _083_ = io_resetMode ? (* src = "CanFifo.scala:46.31" *) 1'h0 : io_wr;
  assign _075_ = io_extendedMode ? (* src = "CanFifo.scala:59.45" *) 6'h10 : 6'h14;
  assign _002_ = _039_ ? (* src = "CanFifo.scala:87.40|CanFifo.scala:88.18" *) 1'h0 : _022_;
  assign _003_ = _050_ ? (* src = "CanFifo.scala:99.65|CanFifo.scala:100.15|CanFifo.scala:48.31" *) _067_ : { 1'h0, fifoCnt };
  assign _004_ = _047_ ? (* src = "CanFifo.scala:97.54|CanFifo.scala:98.13" *) { 1'h0, _066_ } : _003_;
  assign _005_ = _044_ ? (* src = "CanFifo.scala:95.53|CanFifo.scala:96.13" *) _063_ : _004_;
  assign _006_ = io_resetMode ? (* src = "CanFifo.scala:93.22|CanFifo.scala:94.13" *) 8'h00 : _005_;
  assign _007_ = _056_ ? (* src = "CanFifo.scala:108.45|CanFifo.scala:109.15|CanFifo.scala:23.31" *) _069_ : { 1'h0, infoCnt };
  assign _008_ = _053_ ? (* src = "CanFifo.scala:106.44|CanFifo.scala:107.15" *) _068_ : _007_;
  assign _009_ = _051_ ? (* src = "CanFifo.scala:105.50|CanFifo.scala:23.31" *) _008_ : { 1'h0, infoCnt };
  assign _010_ = io_resetMode ? (* src = "CanFifo.scala:103.22|CanFifo.scala:104.13" *) 8'h00 : _009_;
  assign _011_ = _055_ ? (* src = "CanFifo.scala:113.30|CanFifo.scala:114.24|CanFifo.scala:51.42" *) 1'h0 : initializeMemories;
  assign _000_ = _046_ ? (* src = "CanFifo.scala:63.35|CanFifo.scala:64.12|CanFifo.scala:47.30" *) _071_ : lenCnt;
  assign _015_ = reset ? (* src = "CanFifo.scala:23.31|CanFifo.scala:23.31" *) 8'h00 : _010_;
  assign _016_ = reset ? (* src = "CanFifo.scala:45.37|CanFifo.scala:45.37" *) 7'h00 : _018_;
  assign _017_ = reset ? (* src = "CanFifo.scala:48.31|CanFifo.scala:48.31" *) 8'h00 : _006_;
  assign _001_ = _039_ ? (* src = "CanFifo.scala:61.40|CanFifo.scala:62.12" *) 4'h0 : _000_;
  assign _012_ = io_resetMode ? (* src = "CanFifo.scala:69.28|CanFifo.scala:70.19|CanFifo.scala:44.37" *) rdInfoPointer : wrInfoPointer;
  assign _013_ = _059_ ? (* src = "CanFifo.scala:67.60|CanFifo.scala:68.19" *) _080_ : _012_;
  assign _018_ = _060_ ? (* src = "CanFifo.scala:73.38|CanFifo.scala:74.19|CanFifo.scala:45.37" *) _072_ : { 1'h0, rdInfoPointer };
  assign _019_ = _062_ ? (* src = "CanFifo.scala:77.39|CanFifo.scala:78.15|CanFifo.scala:41.33" *) _074_ : rdPointer;
  assign _020_ = _046_ ? (* src = "CanFifo.scala:83.33|CanFifo.scala:84.15|CanFifo.scala:42.33" *) _082_ : wrPointer;
  assign _021_ = io_resetMode ? (* src = "CanFifo.scala:81.22|CanFifo.scala:82.15" *) rdPointer : _020_;
  assign _084_ = ~ io_wr;
  assign _040_ = ~ fifoFull;
  assign _054_ = ~ infoFull;
  assign _061_ = ~ fifoEmpty;
  assign _042_ = ~ io_releaseBuffer;
  assign _052_ = ~ io_infoEmpty;
  assign _058_ = ~ initializeMemories;
  assign _026_ = _056_ | initializeMemories;
  assign _032_ = _056_ | initializeMemories;
  assign _037_ = reset | _011_;
  assign _039_ = io_resetMode | writeLengthInfo;
  assign _059_ = _056_ | initializeMemories;
  assign _022_ = _041_ | latchOverrun;
  assign _057_ = latchOverrun | _041_;
  always @(posedge clock)
    initializeMemories <= _037_;
  always @(posedge clock)
    latchOverrun <= _087_;
  always @(posedge clock)
    fifoCnt <= _017_[6:0];
  always @(posedge clock)
    lenCnt <= _089_;
  always @(posedge clock)
    wrQ <= _091_;
  always @(posedge clock)
    rdInfoPointer <= _016_[5:0];
  always @(posedge clock)
    wrInfoPointer <= _093_;
  always @(posedge clock)
    wrPointer <= _095_;
  always @(posedge clock)
    rdPointer <= _097_;
  always @(posedge clock)
    infoCnt <= _015_[6:0];
  assign _087_ = _088_ ? (* full_case = 32'd1 *) (* src = "CanFifo.scala:50.36" *) 1'h0 : _002_;
  assign _089_ = _090_ ? (* full_case = 32'd1 *) (* src = "CanFifo.scala:47.30" *) 4'h0 : _001_;
  assign _091_ = _092_ ? (* full_case = 32'd1 *) (* src = "CanFifo.scala:46.27" *) 1'h0 : _083_;
  assign _093_ = _094_ ? (* full_case = 32'd1 *) (* src = "CanFifo.scala:44.37" *) 6'h00 : _013_;
  assign _095_ = _096_ ? (* full_case = 32'd1 *) (* src = "CanFifo.scala:42.33" *) 6'h00 : _021_;
  assign _097_ = _098_ ? (* full_case = 32'd1 *) (* src = "CanFifo.scala:41.33" *) 6'h00 : _019_;
  assign _055_ = & wrInfoPointer;
  assign _076_ = { 1'h0, io_addr } - { 1'h0, _075_ };
  assign _065_ = { 1'h0, fifoCnt } - { 1'h0, _064_ };
  assign _068_ = { 1'h0, infoCnt } - 8'h01;
  assign _051_ = writeLengthInfo ^ io_releaseBuffer;
  assign _077_ = _076_[5:0];
  assign _071_ = _070_[3:0];
  assign _080_ = _079_[5:0];
  assign lengthInfo = lengthFifo_lengthInfo_MPORT_data;
  assign _014_ = { 2'h0, lengthInfo };
  assign _074_ = _073_[5:0];
  assign _082_ = _081_[5:0];
  assign _064_ = { 3'h0, lengthInfo };
  assign _066_ = _065_[6:0];
  assign io_dataOut = fifo_io_dataOut_MPORT_data;
  assign io_overrun = overrunInfo_io_overrun_MPORT_data;
  assign io_infoCnt = infoCnt;
  assign \initializeMemories$process$CanFifo_8  = _037_;
  assign \fifoCnt$process$CanFifo_6  = _017_[6:0];
  assign \rdInfoPointer$process$CanFifo_3  = _016_[5:0];
  assign \infoCnt$process$CanFifo  = _015_[6:0];
  assign _088_ = reset;
  assign \latchOverrun$process$CanFifo_7  = _087_;
  assign _090_ = reset;
  assign \lenCnt$process$CanFifo_5  = _089_;
  assign _092_ = reset;
  assign \wrQ$process$CanFifo_4  = _091_;
  assign _094_ = reset;
  assign \wrInfoPointer$process$CanFifo_2  = _093_;
  assign _096_ = reset;
  assign \wrPointer$process$CanFifo_1  = _095_;
  assign _098_ = reset;
  assign \rdPointer$process$CanFifo_0  = _097_;
endmodule

(* cells_not_processed =  1  *)
module CanRegister(clock, reset, io_dataIn, io_dataOut, io_writeEn);
  (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *)
  wire [3:0] _0_;
  wire [3:0] _1_;
  wire _2_;
  input clock;
  (* src = "CanRegister.scala:13.31" *)
  reg [3:0] dataOut;
  (* src = "CanRegister.scala:13.31|CanRegister.scala:13.31" *)
  wire [3:0] \dataOut$process$CanRegister ;
  input [3:0] io_dataIn;
  output [3:0] io_dataOut;
  input io_writeEn;
  input reset;
  assign _0_ = io_writeEn ? (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *) io_dataIn : dataOut;
  always @(posedge clock)
    dataOut <= _1_;
  assign _1_ = _2_ ? (* full_case = 32'd1 *) (* src = "CanRegister.scala:13.31" *) 4'h0 : _0_;
  assign io_dataOut = dataOut;
  assign _2_ = reset;
  assign \dataOut$process$CanRegister  = _1_;
endmodule

(* cells_not_processed =  1  *)
module CanRegisterDoubleReset(clock, reset, io_resetSync, io_dataIn, io_dataOut, io_writeEn);
  (* src = "CanRegisterDoubleReset.scala:17.26|CanRegisterDoubleReset.scala:18.15|CanRegisterDoubleReset.scala:13.31" *)
  wire _0_;
  (* src = "CanRegisterDoubleReset.scala:15.22|CanRegisterDoubleReset.scala:16.13" *)
  wire _1_;
  wire _2_;
  input clock;
  (* src = "CanRegisterDoubleReset.scala:13.31" *)
  reg dataOut;
  (* src = "CanRegisterDoubleReset.scala:13.31|CanRegisterDoubleReset.scala:13.31" *)
  wire \dataOut$process$CanRegisterDoubleReset ;
  input io_dataIn;
  output io_dataOut;
  input io_resetSync;
  input io_writeEn;
  input reset;
  assign _0_ = io_writeEn ? (* src = "CanRegisterDoubleReset.scala:17.26|CanRegisterDoubleReset.scala:18.15|CanRegisterDoubleReset.scala:13.31" *) io_dataIn : dataOut;
  assign _2_ = reset | _1_;
  assign _1_ = io_resetSync | _0_;
  always @(posedge clock)
    dataOut <= _2_;
  assign io_dataOut = dataOut;
  assign \dataOut$process$CanRegisterDoubleReset  = _2_;
endmodule

(* cells_not_processed =  1  *)
module CanRegisterDoubleReset_1(clock, reset, io_resetSync, io_dataIn, io_dataOut, io_writeEn);
  (* src = "CanRegisterDoubleReset.scala:17.26|CanRegisterDoubleReset.scala:18.15|CanRegisterDoubleReset.scala:13.31" *)
  wire _0_;
  (* src = "CanRegisterDoubleReset.scala:15.22|CanRegisterDoubleReset.scala:16.13" *)
  wire _1_;
  wire _2_;
  wire _3_;
  input clock;
  (* src = "CanRegisterDoubleReset.scala:13.31" *)
  reg dataOut;
  (* src = "CanRegisterDoubleReset.scala:13.31|CanRegisterDoubleReset.scala:13.31" *)
  wire \dataOut$process$CanRegisterDoubleReset_1 ;
  input io_dataIn;
  output io_dataOut;
  input io_resetSync;
  input io_writeEn;
  input reset;
  assign _0_ = io_writeEn ? (* src = "CanRegisterDoubleReset.scala:17.26|CanRegisterDoubleReset.scala:18.15|CanRegisterDoubleReset.scala:13.31" *) io_dataIn : dataOut;
  assign _1_ = io_resetSync ? (* src = "CanRegisterDoubleReset.scala:15.22|CanRegisterDoubleReset.scala:16.13" *) 1'h0 : _0_;
  always @(posedge clock)
    dataOut <= _2_;
  assign _2_ = _3_ ? (* full_case = 32'd1 *) (* src = "CanRegisterDoubleReset.scala:13.31" *) 1'h0 : _1_;
  assign io_dataOut = dataOut;
  assign _3_ = reset;
  assign \dataOut$process$CanRegisterDoubleReset_1  = _2_;
endmodule

(* cells_not_processed =  1  *)
module CanRegister_1(clock, reset, io_dataIn, io_dataOut, io_writeEn);
  (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *)
  wire [2:0] _0_;
  wire [2:0] _1_;
  wire _2_;
  input clock;
  (* src = "CanRegister.scala:13.31" *)
  reg [2:0] dataOut;
  (* src = "CanRegister.scala:13.31|CanRegister.scala:13.31" *)
  wire [2:0] \dataOut$process$CanRegister_1 ;
  input [2:0] io_dataIn;
  output [2:0] io_dataOut;
  input io_writeEn;
  input reset;
  assign _0_ = io_writeEn ? (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *) io_dataIn : dataOut;
  always @(posedge clock)
    dataOut <= _1_;
  assign _1_ = _2_ ? (* full_case = 32'd1 *) (* src = "CanRegister.scala:13.31" *) 3'h0 : _0_;
  assign io_dataOut = dataOut;
  assign _2_ = reset;
  assign \dataOut$process$CanRegister_1  = _1_;
endmodule

(* cells_not_processed =  1  *)
module CanRegister_2(clock, reset, io_dataIn, io_dataOut, io_writeEn);
  (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *)
  wire [7:0] _0_;
  wire [7:0] _1_;
  wire _2_;
  input clock;
  (* src = "CanRegister.scala:13.31" *)
  reg [7:0] dataOut;
  (* src = "CanRegister.scala:13.31|CanRegister.scala:13.31" *)
  wire [7:0] \dataOut$process$CanRegister_2 ;
  input [7:0] io_dataIn;
  output [7:0] io_dataOut;
  input io_writeEn;
  input reset;
  assign _0_ = io_writeEn ? (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *) io_dataIn : dataOut;
  always @(posedge clock)
    dataOut <= _1_;
  assign _1_ = _2_ ? (* full_case = 32'd1 *) (* src = "CanRegister.scala:13.31" *) 8'h00 : _0_;
  assign io_dataOut = dataOut;
  assign _2_ = reset;
  assign \dataOut$process$CanRegister_2  = _1_;
endmodule

(* cells_not_processed =  1  *)
module CanRegister_5(clock, reset, io_dataIn, io_dataOut, io_writeEn);
  (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *)
  wire [7:0] _0_;
  wire [7:0] _1_;
  wire _2_;
  input clock;
  (* src = "CanRegister.scala:13.31" *)
  reg [7:0] dataOut;
  (* src = "CanRegister.scala:13.31|CanRegister.scala:13.31" *)
  wire [7:0] \dataOut$process$CanRegister_5 ;
  input [7:0] io_dataIn;
  output [7:0] io_dataOut;
  input io_writeEn;
  input reset;
  assign _0_ = io_writeEn ? (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *) io_dataIn : dataOut;
  always @(posedge clock)
    dataOut <= _1_;
  assign _1_ = _2_ ? (* full_case = 32'd1 *) (* src = "CanRegister.scala:13.31" *) 8'h60 : _0_;
  assign io_dataOut = dataOut;
  assign _2_ = reset;
  assign \dataOut$process$CanRegister_5  = _1_;
endmodule

(* cells_not_processed =  1  *)
module CanRegister_6(clock, reset, io_dataIn, io_dataOut, io_writeEn);
  (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *)
  wire _0_;
  wire _1_;
  wire _2_;
  input clock;
  (* src = "CanRegister.scala:13.31" *)
  reg dataOut;
  (* src = "CanRegister.scala:13.31|CanRegister.scala:13.31" *)
  wire \dataOut$process$CanRegister_6 ;
  input io_dataIn;
  output io_dataOut;
  input io_writeEn;
  input reset;
  assign _0_ = io_writeEn ? (* src = "CanRegister.scala:15.20|CanRegister.scala:16.13|CanRegister.scala:13.31" *) io_dataIn : dataOut;
  always @(posedge clock)
    dataOut <= _1_;
  assign _1_ = _2_ ? (* full_case = 32'd1 *) (* src = "CanRegister.scala:13.31" *) 1'h0 : _0_;
  assign io_dataOut = dataOut;
  assign _2_ = reset;
  assign \dataOut$process$CanRegister_6  = _1_;
endmodule

(* cells_not_processed =  1  *)
module CanRegisters(clock, reset, io_cs, io_writeEn, io_addr, io_dataIn, io_dataOut, io_irqN, io_samplePoint, io_transmitting, io_setResetMode, io_nodeBusOff, io_errorStatus, io_rxErrorCount, io_txErrorCount, io_transmitStatus, io_receiveStatus, io_txSuccessful, io_needToTx, io_overrun, io_infoEmpty
, io_setBusErrorIrq, io_setArbitrationLostIrq, io_arbitrationLostCapture, io_nodeErrorPassive, io_nodeErrorActive, io_rxMessageCounter, io_resetMode, io_listenOnlyMode, io_acceptanceFilterMode, io_selfTestMode, io_clearDataOverrun, io_releaseBuffer, io_abortTx, io_txRequest, io_selfRxRequest, io_singleShotTransmission, io_txState, io_txStateQ, io_overloadFrame, io_readArbitrationLostCaptureReg, io_readErrorCodeCaptureReg
, io_errorCaptureCode, io_baudRatePrescaler, io_syncJumpWidth, io_timeSegment1, io_timeSegment2, io_tripleSampling, io_errorWarningLimit, io_writeEnReceiveErrorCounter, io_writeEnTransmitErrorCounter, io_extendedMode, io_clkout, io_acceptanceCode_0, io_acceptanceCode_1, io_acceptanceCode_2, io_acceptanceCode_3, io_acceptanceMask_0, io_acceptanceMask_1, io_acceptanceMask_2, io_acceptanceMask_3, io_txData_0, io_txData_1
, io_txData_2, io_txData_3, io_txData_4, io_txData_5, io_txData_6, io_txData_7, io_txData_8, io_txData_9, io_txData_10, io_txData_11, io_txData_12);
  (* src = "CanRegisters.scala:182.43|CanRegisters.scala:183.19|CanRegisters.scala:102.36" *)
  wire _000_;
  (* src = "CanRegisters.scala:180.34|CanRegisters.scala:181.19" *)
  wire _001_;
  (* src = "CanRegisters.scala:235.28|CanRegisters.scala:236.25|CanRegisters.scala:112.42" *)
  wire _002_;
  (* src = "CanRegisters.scala:232.41|CanRegisters.scala:233.25" *)
  wire _003_;
  (* src = "CanRegisters.scala:271.33|CanRegisters.scala:272.15|CanRegisters.scala:276.15" *)
  wire [2:0] _004_;
  (* src = "CanRegisters.scala:271.33|CanRegisters.scala:273.15|CanRegisters.scala:269.33" *)
  wire _005_;
  (* src = "CanRegisters.scala:358.41|CanRegisters.scala:359.20|CanRegisters.scala:348.38" *)
  wire _006_;
  (* src = "CanRegisters.scala:356.51|CanRegisters.scala:357.20" *)
  wire _007_;
  (* src = "CanRegisters.scala:364.77|CanRegisters.scala:365.17|CanRegisters.scala:349.35" *)
  wire _008_;
  (* src = "CanRegisters.scala:362.35|CanRegisters.scala:363.17" *)
  wire _009_;
  (* src = "CanRegisters.scala:370.48|CanRegisters.scala:371.16|CanRegisters.scala:350.34" *)
  wire _010_;
  (* src = "CanRegisters.scala:194.42|CanRegisters.scala:195.28|CanRegisters.scala:104.45" *)
  wire _011_;
  (* src = "CanRegisters.scala:368.56|CanRegisters.scala:369.16" *)
  wire _012_;
  (* src = "CanRegisters.scala:376.26|CanRegisters.scala:377.14|CanRegisters.scala:351.32" *)
  wire _013_;
  (* src = "CanRegisters.scala:374.95|CanRegisters.scala:375.14" *)
  wire _014_;
  (* src = "CanRegisters.scala:382.41|CanRegisters.scala:383.17|CanRegisters.scala:352.35" *)
  wire _015_;
  (* src = "CanRegisters.scala:380.43|CanRegisters.scala:381.17" *)
  wire _016_;
  (* src = "CanRegisters.scala:388.41|CanRegisters.scala:389.24|CanRegisters.scala:353.42" *)
  wire _017_;
  (* src = "CanRegisters.scala:386.57|CanRegisters.scala:387.24" *)
  wire _018_;
  (* src = "CanRegisters.scala:394.41|CanRegisters.scala:395.21|CanRegisters.scala:354.39" *)
  wire _019_;
  (* src = "CanRegisters.scala:392.140|CanRegisters.scala:393.21" *)
  wire _020_;
  (* src = "CanRegisters.scala:403.19|CanRegisters.scala:404.10|CanRegisters.scala:100.27" *)
  wire _021_;
  (* src = "CanRegisters.scala:191.52|CanRegisters.scala:192.28" *)
  wire _022_;
  (* src = "CanRegisters.scala:401.39|CanRegisters.scala:402.10" *)
  wire _023_;
  (* src = "CanRegisters.scala:214.43|CanRegisters.scala:215.26|CanRegisters.scala:110.43" *)
  wire _024_;
  (* src = "CanRegisters.scala:212.22|CanRegisters.scala:213.26" *)
  wire _025_;
  (* src = "CanRegisters.scala:221.27|CanRegisters.scala:222.26|CanRegisters.scala:109.43" *)
  wire _026_;
  (* src = "CanRegisters.scala:218.57|CanRegisters.scala:219.26" *)
  wire _027_;
  (* src = "CanRegisters.scala:228.49|CanRegisters.scala:229.19|CanRegisters.scala:108.36" *)
  wire _028_;
  (* src = "CanRegisters.scala:225.32|CanRegisters.scala:226.19" *)
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire [1:0] _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire [2:0] _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire [3:0] _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire [1:0] _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire [1:0] _064_;
  wire [1:0] _065_;
  wire [1:0] _066_;
  wire [1:0] _067_;
  wire [3:0] _068_;
  wire [1:0] _069_;
  wire [1:0] _070_;
  wire [1:0] _071_;
  wire [1:0] _072_;
  wire [1:0] _073_;
  wire [1:0] _074_;
  wire [3:0] _075_;
  wire [1:0] _076_;
  wire [1:0] _077_;
  wire [1:0] _078_;
  wire [1:0] _079_;
  wire [1:0] _080_;
  wire [3:0] _081_;
  wire [1:0] _082_;
  wire [1:0] _083_;
  wire [1:0] _084_;
  wire [3:0] _085_;
  wire [3:0] _086_;
  wire [3:0] _087_;
  wire [3:0] _088_;
  wire [3:0] _089_;
  wire [6:0] _090_;
  wire [6:0] _091_;
  wire [6:0] _092_;
  wire [1:0] _093_;
  wire [1:0] _094_;
  wire [1:0] _095_;
  wire [1:0] _096_;
  wire [3:0] _097_;
  wire [1:0] _098_;
  wire [1:0] _099_;
  wire [1:0] _100_;
  wire [1:0] _101_;
  wire [1:0] _102_;
  wire [3:0] _103_;
  wire [3:0] _104_;
  wire [1:0] _105_;
  wire [1:0] _106_;
  wire [1:0] _107_;
  wire [1:0] _108_;
  wire [1:0] _109_;
  wire [3:0] _110_;
  wire [1:0] _111_;
  wire [1:0] _112_;
  wire [1:0] _113_;
  wire [1:0] _114_;
  wire [1:0] _115_;
  wire [1:0] _116_;
  wire [3:0] _117_;
  wire [1:0] _118_;
  wire [1:0] _119_;
  wire [1:0] _120_;
  wire [1:0] _121_;
  wire [1:0] _122_;
  wire [3:0] _123_;
  wire [1:0] _124_;
  wire [1:0] _125_;
  wire [1:0] _126_;
  wire [6:0] _127_;
  wire [6:0] _128_;
  wire [6:0] _129_;
  wire _130_;
  wire _131_;
  wire [3:0] _132_;
  wire _133_;
  wire [2:0] _134_;
  wire _135_;
  wire _136_;
  wire [1:0] _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire [1:0] _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  (* src = "CanRegisters.scala:180.21" *)
  wire _159_;
  (* src = "CanRegisters.scala:180.19" *)
  wire _160_;
  (* src = "CanRegisters.scala:218.27" *)
  wire _161_;
  (* src = "CanRegisters.scala:218.24" *)
  wire _162_;
  (* src = "CanRegisters.scala:218.43" *)
  wire _163_;
  (* src = "CanRegisters.scala:225.21" *)
  wire _164_;
  (* src = "CanRegisters.scala:225.19" *)
  wire _165_;
  (* src = "CanRegisters.scala:228.26" *)
  wire _166_;
  (* src = "CanRegisters.scala:232.21" *)
  wire _167_;
  (* src = "CanRegisters.scala:235.13" *)
  wire _168_;
  (* src = "CanRegisters.scala:271.18" *)
  wire _169_;
  (* src = "CanRegisters.scala:182.15" *)
  wire _170_;
  (* src = "CanRegisters.scala:356.31" *)
  wire _171_;
  (* src = "CanRegisters.scala:358.27" *)
  wire _172_;
  (* src = "CanRegisters.scala:364.37" *)
  wire _173_;
  (* src = "CanRegisters.scala:364.35" *)
  wire _174_;
  (* src = "CanRegisters.scala:364.60" *)
  wire _175_;
  (* src = "CanRegisters.scala:182.28" *)
  wire _176_;
  (* src = "CanRegisters.scala:368.27" *)
  wire _177_;
  (* src = "CanRegisters.scala:368.24" *)
  wire _178_;
  (* src = "CanRegisters.scala:368.40" *)
  wire _179_;
  (* src = "CanRegisters.scala:374.25" *)
  wire _180_;
  (* src = "CanRegisters.scala:374.58" *)
  wire _181_;
  (* src = "CanRegisters.scala:374.41" *)
  wire _182_;
  (* src = "CanRegisters.scala:374.74" *)
  wire _183_;
  (* src = "CanRegisters.scala:380.26" *)
  wire _184_;
  (* src = "CanRegisters.scala:191.21" *)
  wire _185_;
  (* src = "CanRegisters.scala:386.33" *)
  wire _186_;
  (* src = "CanRegisters.scala:392.32" *)
  wire _187_;
  (* src = "CanRegisters.scala:392.29" *)
  wire _188_;
  (* src = "CanRegisters.scala:392.55" *)
  wire _189_;
  (* src = "CanRegisters.scala:392.77" *)
  wire _190_;
  (* src = "CanRegisters.scala:392.97" *)
  wire _191_;
  (* src = "CanRegisters.scala:392.52" *)
  wire _192_;
  (* src = "CanRegisters.scala:392.119" *)
  wire _193_;
  (* src = "CanRegisters.scala:191.34" *)
  wire _194_;
  (* src = "CanRegisters.scala:401.19" *)
  wire _195_;
  (* src = "CanRegisters.scala:214.29" *)
  wire _196_;
  (* src = "CanRegisters.scala:214.27" *)
  wire _197_;
  (* src = "CanRegisters.scala:276.28" *)
  wire [3:0] _198_;
  (* src = "CanRegisters.scala:276.28" *)
  wire [2:0] _199_;
  (* src = "CanRegisters.scala:266.33" *)
  wire _200_;
  (* src = "CanRegisters.scala:273.18" *)
  wire _201_;
  (* src = "CanRegisters.scala:174.53" *)
  wire _202_;
  (* src = "CanRegisters.scala:175.89" *)
  wire _203_;
  (* src = "CanRegisters.scala:175.87" *)
  wire _204_;
  (* src = "CanRegisters.scala:175.73" *)
  wire _205_;
  (* src = "CanRegisters.scala:175.57" *)
  wire _206_;
  (* src = "CanRegisters.scala:176.53" *)
  wire _207_;
  (* src = "CanRegisters.scala:178.53" *)
  wire _208_;
  (* src = "CanRegisters.scala:189.30" *)
  wire _209_;
  (* src = "CanRegisters.scala:171.55" *)
  wire _210_;
  (* src = "CanRegisters.scala:279.50" *)
  wire _211_;
  (* src = "CanRegisters.scala:279.66" *)
  wire _212_;
  (* src = "CanRegisters.scala:282.28" *)
  wire _213_;
  (* src = "CanRegisters.scala:285.27" *)
  wire _214_;
  (* src = "CanRegisters.scala:298.22" *)
  wire [4:0] _215_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _216_;
  (* src = "Mux.scala:80.60" *)
  wire _217_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _218_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _219_;
  (* src = "Mux.scala:80.60" *)
  wire _220_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _221_;
  (* src = "Mux.scala:80.60" *)
  wire _222_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _223_;
  (* src = "Mux.scala:80.60" *)
  wire _224_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _225_;
  (* src = "Mux.scala:80.60" *)
  wire _226_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _227_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _228_;
  (* src = "Mux.scala:80.60" *)
  wire _229_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _230_;
  (* src = "Mux.scala:80.60" *)
  wire _231_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _232_;
  (* src = "Mux.scala:80.60" *)
  wire _233_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _234_;
  (* src = "Mux.scala:80.60" *)
  wire _235_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _236_;
  (* src = "Mux.scala:80.60" *)
  wire _237_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _238_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _239_;
  (* src = "Mux.scala:80.60" *)
  wire _240_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _241_;
  (* src = "Mux.scala:80.60" *)
  wire _242_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _243_;
  (* src = "Mux.scala:80.60" *)
  wire _244_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _245_;
  (* src = "Mux.scala:80.60" *)
  wire _246_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _247_;
  (* src = "Mux.scala:80.60" *)
  wire _248_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _249_;
  (* src = "Mux.scala:80.60" *)
  wire _250_;
  (* src = "Mux.scala:80.60" *)
  wire _251_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _252_;
  (* src = "Mux.scala:80.60" *)
  wire _253_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _254_;
  (* src = "Mux.scala:80.60" *)
  wire _255_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _256_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _257_;
  (* src = "CanRegisters.scala:325.35" *)
  wire [3:0] _258_;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] _259_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _260_;
  (* src = "CanRegisters.scala:326.17" *)
  wire [7:0] _261_;
  (* src = "CanRegisters.scala:327.17" *)
  wire [7:0] _262_;
  (* src = "CanRegisters.scala:328.17" *)
  wire [7:0] _263_;
  (* src = "CanRegisters.scala:329.17" *)
  wire [7:0] _264_;
  (* src = "CanRegisters.scala:330.18" *)
  wire [7:0] _265_;
  (* src = "CanRegisters.scala:331.18" *)
  wire [7:0] _266_;
  (* src = "CanRegisters.scala:332.18" *)
  wire [7:0] _267_;
  (* src = "CanRegisters.scala:333.18" *)
  wire [7:0] _268_;
  (* src = "CanRegisters.scala:334.18" *)
  wire [7:0] _269_;
  (* src = "CanRegisters.scala:335.18" *)
  wire [7:0] _270_;
  (* src = "Mux.scala:80.60" *)
  wire _271_;
  (* src = "CanRegisters.scala:336.18" *)
  wire [7:0] _272_;
  (* src = "CanRegisters.scala:337.18" *)
  wire [7:0] _273_;
  (* src = "CanRegisters.scala:338.18" *)
  wire [7:0] _274_;
  (* src = "CanRegisters.scala:339.18" *)
  wire [7:0] _275_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _276_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _277_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _278_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _279_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _280_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _281_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _282_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _283_;
  (* src = "Mux.scala:80.60" *)
  wire _284_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _285_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _286_;
  (* src = "Mux.scala:80.60" *)
  wire _287_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _288_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _289_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _290_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _291_;
  (* src = "Mux.scala:80.60" *)
  wire _292_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _293_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _294_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _295_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _296_;
  (* src = "Mux.scala:80.60" *)
  wire _297_;
  (* src = "Mux.scala:80.57" *)
  wire [7:0] _298_;
  (* src = "CanRegisters.scala:169.49" *)
  wire _299_;
  (* src = "CanRegisters.scala:200.69" *)
  wire _300_;
  (* src = "CanRegisters.scala:134.44" *)
  wire _301_;
  (* src = "CanRegisters.scala:134.73" *)
  wire _302_;
  (* src = "CanRegisters.scala:135.67" *)
  wire _303_;
  (* src = "CanRegisters.scala:170.47" *)
  wire _304_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _305_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _306_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _307_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _308_;
  (* src = "CanRegisters.scala:133.42" *)
  wire _309_;
  (* src = "CanRegisters.scala:132.29" *)
  wire _310_;
  (* src = "CanRegisters.scala:93.28" *)
  wire _311_;
  (* src = "CanRegisters.scala:93.57" *)
  wire _312_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _313_;
  (* src = "CanRegisters.scala:93.107" *)
  wire _314_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _315_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _316_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _317_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _318_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _319_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _320_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _321_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _322_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _323_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _324_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _325_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _326_;
  (* src = "CanRegisters.scala:93.57" *)
  wire _327_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _328_;
  (* src = "CanRegisters.scala:93.107" *)
  wire _329_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _330_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _331_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _332_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _333_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _334_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _335_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _336_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _337_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _338_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _339_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _340_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _341_;
  (* src = "CanRegisters.scala:97.35" *)
  wire _342_;
  (* src = "CanRegisters.scala:97.24" *)
  wire _343_;
  (* src = "CanRegisters.scala:97.35" *)
  wire _344_;
  (* src = "CanRegisters.scala:97.24" *)
  wire _345_;
  (* src = "CanRegisters.scala:97.35" *)
  wire _346_;
  (* src = "CanRegisters.scala:97.35" *)
  wire _347_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _348_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _349_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _350_;
  (* src = "CanRegisters.scala:97.11" *)
  wire _351_;
  (* src = "CanRegisters.scala:97.35" *)
  wire _352_;
  (* src = "CanRegisters.scala:93.57" *)
  wire _353_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _354_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _355_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _356_;
  (* src = "CanRegisters.scala:150.61" *)
  wire _357_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _358_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _359_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _360_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _361_;
  (* src = "CanRegisters.scala:152.48" *)
  wire _362_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _363_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _364_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _365_;
  (* src = "CanRegisters.scala:152.48" *)
  wire _366_;
  (* src = "CanRegisters.scala:89.35" *)
  wire _367_;
  (* src = "CanRegisters.scala:89.24" *)
  wire _368_;
  (* src = "CanRegisters.scala:89.59" *)
  wire _369_;
  (* src = "CanRegisters.scala:152.48" *)
  wire _370_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _371_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _372_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _373_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _374_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _375_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _376_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _377_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _378_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _379_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _380_;
  (* src = "CanRegisters.scala:93.57" *)
  wire _381_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _382_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _383_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _384_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _385_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _386_;
  (* src = "CanRegisters.scala:93.57" *)
  wire _387_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _388_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _389_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _390_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _391_;
  (* src = "CanRegisters.scala:93.57" *)
  wire _392_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _393_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _394_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _395_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _396_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _397_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _398_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _399_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _400_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _401_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _402_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _403_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _404_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _405_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _406_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _407_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _408_;
  (* src = "CanRegisters.scala:93.107" *)
  wire _409_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _410_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _411_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _412_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _413_;
  (* src = "CanRegisters.scala:93.46" *)
  wire _414_;
  (* src = "CanRegisters.scala:93.107" *)
  wire _415_;
  (* src = "CanRegisters.scala:93.96" *)
  wire _416_;
  (* src = "CanRegisters.scala:93.78" *)
  wire _417_;
  (* src = "CanRegisters.scala:93.24" *)
  wire _418_;
  (* src = "CanRegisters.scala:150.58" *)
  wire _419_;
  wire _420_;
  wire _421_;
  wire _422_;
  wire _423_;
  wire _424_;
  wire _425_;
  wire _426_;
  wire _427_;
  wire _428_;
  wire _429_;
  wire _430_;
  wire _431_;
  wire _432_;
  wire _433_;
  wire _434_;
  wire _435_;
  wire [2:0] _436_;
  wire _437_;
  wire _438_;
  wire _439_;
  wire _440_;
  wire _441_;
  wire _442_;
  wire _443_;
  wire _444_;
  wire _445_;
  wire _446_;
  wire _447_;
  (* src = "CanRegisters.scala:353.42" *)
  reg arbitrationLostIrq;
  (* src = "CanRegisters.scala:353.42|CanRegisters.scala:353.42" *)
  wire \arbitrationLostIrq$process$CanRegisters_16 ;
  (* src = "CanRegisters.scala:241.45" *)
  wire arbitrationLostIrqEn;
  (* src = "CanRegisters.scala:352.35" *)
  reg busErrorIrq;
  (* src = "CanRegisters.scala:352.35|CanRegisters.scala:352.35" *)
  wire \busErrorIrq$process$CanRegisters_15 ;
  (* src = "CanRegisters.scala:240.38" *)
  wire busErrorIrqEn;
  wire [7:0] busTiming0_m_io_dataOut;
  wire [7:0] busTiming1_m_io_dataOut;
  wire [2:0] cd_m_io_dataOut;
  (* src = "CanRegisters.scala:268.33" *)
  reg [2:0] clkoutCnt;
  (* src = "CanRegisters.scala:268.33|CanRegisters.scala:268.33" *)
  wire [2:0] \clkoutCnt$process$CanRegisters_13 ;
  (* src = "CanRegisters.scala:266.29" *)
  wire [2:0] clkoutDiv;
  (* src = "CanRegisters.scala:269.33" *)
  reg clkoutTmp;
  (* src = "CanRegisters.scala:269.33|CanRegisters.scala:269.33" *)
  wire \clkoutTmp$process$CanRegisters_14 ;
  input clock;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] clockDivider;
  (* src = "CanRegisters.scala:264.79" *)
  wire clockOff;
  (* src = "CanRegisters.scala:264.79" *)
  wire clockOff_m_io_dataOut;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:174.14" *)
  wire command_0;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:174.14" *)
  wire command_0_m_io_dataOut;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:175.14" *)
  wire command_1;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:175.14" *)
  wire command_1_m_io_dataOut;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:176.14" *)
  wire command_2;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:176.14" *)
  wire command_2_m_io_dataOut;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:177.14" *)
  wire command_3;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:177.14" *)
  wire command_3_m_io_dataOut;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:178.14" *)
  wire command_4;
  (* src = "CanRegisters.scala:173.32|CanRegisters.scala:178.14" *)
  wire command_4_m_io_dataOut;
  (* src = "CanRegisters.scala:348.38" *)
  reg dataOverrunIrq;
  (* src = "CanRegisters.scala:348.38|CanRegisters.scala:348.38" *)
  wire \dataOverrunIrq$process$CanRegisters_18 ;
  (* src = "CanRegisters.scala:343.26" *)
  wire dataOverrunIrqEn;
  (* src = "CanRegisters.scala:243.44" *)
  wire dataOverrunIrqEnExt;
  (* src = "CanRegisters.scala:351.32" *)
  reg errorIrq;
  (* src = "CanRegisters.scala:351.32|CanRegisters.scala:351.32" *)
  wire \errorIrq$process$CanRegisters_19 ;
  (* src = "CanRegisters.scala:165.40" *)
  wire errorIrqEnBasic;
  (* src = "CanRegisters.scala:354.39" *)
  reg errorPassiveIrq;
  (* src = "CanRegisters.scala:354.39|CanRegisters.scala:354.39" *)
  wire \errorPassiveIrq$process$CanRegisters_17 ;
  (* src = "CanRegisters.scala:242.42" *)
  wire errorPassiveIrqEn;
  (* src = "CanRegisters.scala:113.35" *)
  reg errorStatusQ;
  (* src = "CanRegisters.scala:113.35" *)
  wire \errorStatusQ$process$CanRegisters_9 ;
  (* src = "CanRegisters.scala:344.27" *)
  wire errorWarningIrqEn;
  (* src = "CanRegisters.scala:244.45" *)
  wire errorWarningIrqEnExt;
  output io_abortTx;
  output [7:0] io_acceptanceCode_0;
  (* src = "CanRegisters.scala:289.26" *)
  wire [7:0] io_acceptanceCode_0_m_io_dataOut;
  output [7:0] io_acceptanceCode_1;
  (* src = "CanRegisters.scala:289.26" *)
  wire [7:0] io_acceptanceCode_1_m_io_dataOut;
  output [7:0] io_acceptanceCode_2;
  (* src = "CanRegisters.scala:289.26" *)
  wire [7:0] io_acceptanceCode_2_m_io_dataOut;
  output [7:0] io_acceptanceCode_3;
  (* src = "CanRegisters.scala:289.26" *)
  wire [7:0] io_acceptanceCode_3_m_io_dataOut;
  output io_acceptanceFilterMode;
  output [7:0] io_acceptanceMask_0;
  (* src = "CanRegisters.scala:290.26" *)
  wire [7:0] io_acceptanceMask_0_m_io_dataOut;
  output [7:0] io_acceptanceMask_1;
  (* src = "CanRegisters.scala:290.26" *)
  wire [7:0] io_acceptanceMask_1_m_io_dataOut;
  output [7:0] io_acceptanceMask_2;
  (* src = "CanRegisters.scala:290.26" *)
  wire [7:0] io_acceptanceMask_2_m_io_dataOut;
  output [7:0] io_acceptanceMask_3;
  (* src = "CanRegisters.scala:290.26" *)
  wire [7:0] io_acceptanceMask_3_m_io_dataOut;
  input [7:0] io_addr;
  input [4:0] io_arbitrationLostCapture;
  output [5:0] io_baudRatePrescaler;
  output io_clearDataOverrun;
  output io_clkout;
  input io_cs;
  input [7:0] io_dataIn;
  output [7:0] io_dataOut;
  input [7:0] io_errorCaptureCode;
  input io_errorStatus;
  output [7:0] io_errorWarningLimit;
  (* src = "CanRegisters.scala:261.24" *)
  wire [7:0] io_errorWarningLimit_m_io_dataOut;
  output io_extendedMode;
  (* src = "CanRegisters.scala:263.76" *)
  wire io_extendedMode_m_io_dataOut;
  input io_infoEmpty;
  output io_irqN;
  output io_listenOnlyMode;
  input io_needToTx;
  input io_nodeBusOff;
  input io_nodeErrorActive;
  input io_nodeErrorPassive;
  input io_overloadFrame;
  input io_overrun;
  output io_readArbitrationLostCaptureReg;
  output io_readErrorCodeCaptureReg;
  input io_receiveStatus;
  output io_releaseBuffer;
  output io_resetMode;
  input [7:0] io_rxErrorCount;
  input [6:0] io_rxMessageCounter;
  input io_samplePoint;
  output io_selfRxRequest;
  output io_selfTestMode;
  input io_setArbitrationLostIrq;
  input io_setBusErrorIrq;
  input io_setResetMode;
  output io_singleShotTransmission;
  output [1:0] io_syncJumpWidth;
  output [3:0] io_timeSegment1;
  output [2:0] io_timeSegment2;
  input io_transmitStatus;
  input io_transmitting;
  output io_tripleSampling;
  output [7:0] io_txData_0;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_0_m_io_dataOut;
  output [7:0] io_txData_1;
  output [7:0] io_txData_10;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_10_m_io_dataOut;
  output [7:0] io_txData_11;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_11_m_io_dataOut;
  output [7:0] io_txData_12;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_12_m_io_dataOut;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_1_m_io_dataOut;
  output [7:0] io_txData_2;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_2_m_io_dataOut;
  output [7:0] io_txData_3;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_3_m_io_dataOut;
  output [7:0] io_txData_4;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_4_m_io_dataOut;
  output [7:0] io_txData_5;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_5_m_io_dataOut;
  output [7:0] io_txData_6;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_6_m_io_dataOut;
  output [7:0] io_txData_7;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_7_m_io_dataOut;
  output [7:0] io_txData_8;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_8_m_io_dataOut;
  output [7:0] io_txData_9;
  (* src = "CanRegisters.scala:294.18" *)
  wire [7:0] io_txData_9_m_io_dataOut;
  input [7:0] io_txErrorCount;
  output io_txRequest;
  input io_txState;
  input io_txStateQ;
  input io_txSuccessful;
  input io_writeEn;
  output io_writeEnReceiveErrorCounter;
  output io_writeEnTransmitErrorCounter;
  (* src = "CanRegisters.scala:399.20" *)
  wire irq;
  (* src = "CanRegisters.scala:239.29|CanRegisters.scala:248.12" *)
  wire [7:0] irqEnExt;
  (* src = "CanRegisters.scala:239.29|CanRegisters.scala:248.12" *)
  wire [7:0] irqEnExt_m_io_dataOut;
  (* src = "CanRegisters.scala:100.27" *)
  reg irqN;
  (* src = "CanRegisters.scala:100.27|CanRegisters.scala:100.27" *)
  wire \irqN$process$CanRegisters ;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] irqReg;
  (* src = "CanRegisters.scala:160.93" *)
  wire mode;
  wire [3:0] modeBasic_m_io_dataOut;
  wire [2:0] modeExt_m_io_dataOut;
  (* src = "CanRegisters.scala:160.93" *)
  wire mode_m_io_dataOut;
  (* src = "CanRegisters.scala:114.34" *)
  reg nodeBusOffQ;
  (* src = "CanRegisters.scala:114.34" *)
  wire \nodeBusOffQ$process$CanRegisters_10 ;
  (* src = "CanRegisters.scala:115.40" *)
  reg nodeErrorPassiveQ;
  (* src = "CanRegisters.scala:115.40" *)
  wire \nodeErrorPassiveQ$process$CanRegisters_11 ;
  (* src = "CanRegisters.scala:198.38" *)
  reg overloadFrameQ;
  (* src = "CanRegisters.scala:198.38|CanRegisters.scala:198.38|CanRegisters.scala:198.38" *)
  wire \overloadFrameQ$process$CanRegisters_12 ;
  (* src = "CanRegisters.scala:166.42" *)
  wire overrunIrqEnBasic;
  (* src = "CanRegisters.scala:107.31" *)
  reg overrunQ;
  (* src = "CanRegisters.scala:107.31" *)
  wire \overrunQ$process$CanRegisters_3 ;
  (* src = "CanRegisters.scala:108.36" *)
  reg overrunStatus;
  (* src = "CanRegisters.scala:108.36|CanRegisters.scala:108.36" *)
  wire \overrunStatus$process$CanRegisters_4 ;
  (* src = "CanRegisters.scala:132.26" *)
  wire read;
  (* src = "CanRegisters.scala:133.31" *)
  wire readIrqReg;
  (* src = "CanRegisters.scala:112.42" *)
  reg receiveBufferStatus;
  (* src = "CanRegisters.scala:112.42|CanRegisters.scala:112.42" *)
  wire \receiveBufferStatus$process$CanRegisters_8 ;
  (* src = "CanRegisters.scala:350.34" *)
  reg receiveIrq;
  (* src = "CanRegisters.scala:350.34|CanRegisters.scala:350.34" *)
  wire \receiveIrq$process$CanRegisters_21 ;
  (* src = "CanRegisters.scala:346.22" *)
  wire receiveIrqEn;
  (* src = "CanRegisters.scala:163.42" *)
  wire receiveIrqEnBasic;
  (* src = "CanRegisters.scala:246.40" *)
  wire receiveIrqEnExt;
  input reset;
  (* src = "CanRegisters.scala:102.36" *)
  reg selfRxRequest;
  (* src = "CanRegisters.scala:102.36|CanRegisters.scala:102.36" *)
  wire \selfRxRequest$process$CanRegisters_0 ;
  (* src = "CanRegisters.scala:104.45" *)
  reg singleShotTransmission;
  (* src = "CanRegisters.scala:104.45|CanRegisters.scala:104.45" *)
  wire \singleShotTransmission$process$CanRegisters_1 ;
  (* src = "Cat.scala:30.58" *)
  wire [7:0] status;
  (* src = "CanRegisters.scala:109.43" *)
  reg transmissionComplete;
  (* src = "CanRegisters.scala:109.43|CanRegisters.scala:109.43" *)
  wire \transmissionComplete$process$CanRegisters_5 ;
  (* src = "CanRegisters.scala:110.43" *)
  reg transmitBufferStatus;
  (* src = "CanRegisters.scala:110.43|CanRegisters.scala:110.43" *)
  wire \transmitBufferStatus$process$CanRegisters_6 ;
  (* src = "CanRegisters.scala:111.44" *)
  reg transmitBufferStatusQ;
  (* src = "CanRegisters.scala:111.44" *)
  wire \transmitBufferStatusQ$process$CanRegisters_7 ;
  (* src = "CanRegisters.scala:349.35" *)
  reg transmitIrq;
  (* src = "CanRegisters.scala:349.35|CanRegisters.scala:349.35" *)
  wire \transmitIrq$process$CanRegisters_20 ;
  (* src = "CanRegisters.scala:345.23" *)
  wire transmitIrqEn;
  (* src = "CanRegisters.scala:164.43" *)
  wire transmitIrqEnBasic;
  (* src = "CanRegisters.scala:245.41" *)
  wire transmitIrqEnExt;
  (* src = "CanRegisters.scala:106.36" *)
  reg txSuccessfulQ;
  (* src = "CanRegisters.scala:106.36" *)
  wire \txSuccessfulQ$process$CanRegisters_2 ;
  (* src = "CanRegisters.scala:97.24" *)
  wire writeEnClockDivLow;
  (* src = "CanRegisters.scala:97.24" *)
  wire writeEnMode;
  assign _198_ = { 1'h0, clkoutCnt } + 4'h1;
  assign _351_ = io_cs & io_writeEn;
  assign writeEnMode = _351_ & _352_;
  assign _343_ = _351_ & _342_;
  assign _328_ = _311_ & _327_;
  assign _193_ = _192_ & errorPassiveIrqEn;
  assign io_listenOnlyMode = io_extendedMode & _299_;
  assign io_acceptanceFilterMode = io_extendedMode & _210_;
  assign io_selfTestMode = io_extendedMode & _304_;
  assign io_abortTx = command_1 & _209_;
  assign io_readArbitrationLostCaptureReg = _301_ & _302_;
  assign io_readErrorCodeCaptureReg = _301_ & _303_;
  assign io_writeEnReceiveErrorCounter = _306_ & io_resetMode;
  assign io_writeEnTransmitErrorCounter = _308_ & io_resetMode;
  assign _131_ = _351_ & _352_;
  assign _330_ = io_extendedMode & _329_;
  assign _133_ = _351_ & _352_;
  assign _135_ = writeEnMode & io_resetMode;
  assign _139_ = _351_ & _347_;
  assign _142_ = _351_ & _347_;
  assign _145_ = _351_ & _347_;
  assign _149_ = _351_ & _347_;
  assign _152_ = _351_ & _347_;
  assign _153_ = io_overloadFrame & _300_;
  assign _155_ = _351_ & _347_;
  assign _156_ = _350_ & io_extendedMode;
  assign _332_ = _351_ & _331_;
  assign _157_ = _343_ & io_resetMode;
  assign _158_ = _345_ & io_resetMode;
  assign _034_ = _349_ & io_resetMode;
  assign _036_ = writeEnClockDivLow & io_resetMode;
  assign _038_ = writeEnClockDivLow & io_resetMode;
  assign _040_ = _351_ & _346_;
  assign _041_ = _317_ & io_resetMode;
  assign _042_ = _332_ & io_resetMode;
  assign _043_ = _320_ & io_resetMode;
  assign _045_ = _335_ & io_resetMode;
  assign _319_ = _351_ & _318_;
  assign _046_ = _323_ & io_resetMode;
  assign _047_ = _338_ & io_resetMode;
  assign _048_ = _326_ & io_resetMode;
  assign _049_ = _341_ & io_resetMode;
  assign _050_ = _358_ & transmitBufferStatus;
  assign _051_ = _375_ & transmitBufferStatus;
  assign _052_ = _380_ & transmitBufferStatus;
  assign _053_ = _386_ & transmitBufferStatus;
  assign _054_ = _391_ & transmitBufferStatus;
  assign _056_ = _397_ & transmitBufferStatus;
  assign _320_ = _319_ & io_extendedMode;
  assign _057_ = _402_ & transmitBufferStatus;
  assign _058_ = _407_ & transmitBufferStatus;
  assign _059_ = _413_ & transmitBufferStatus;
  assign _060_ = _419_ & transmitBufferStatus;
  assign _061_ = _362_ & transmitBufferStatus;
  assign _062_ = _366_ & transmitBufferStatus;
  assign _063_ = _370_ & transmitBufferStatus;
  assign _334_ = _351_ & _333_;
  assign _335_ = _334_ & io_extendedMode;
  assign _322_ = _351_ & _321_;
  assign _323_ = _322_ & io_extendedMode;
  assign _337_ = _351_ & _336_;
  assign _345_ = _351_ & _344_;
  assign _338_ = _337_ & io_extendedMode;
  assign _325_ = _351_ & _324_;
  assign _326_ = _325_ & io_extendedMode;
  assign _340_ = _351_ & _339_;
  assign _341_ = _340_ & io_extendedMode;
  assign _354_ = _311_ & _353_;
  assign _356_ = _351_ & _355_;
  assign _358_ = _356_ & _357_;
  assign _371_ = _311_ & _302_;
  assign _372_ = io_extendedMode & _318_;
  assign writeEnClockDivLow = _351_ & _346_;
  assign _374_ = _351_ & _373_;
  assign _375_ = _374_ & _357_;
  assign _376_ = _311_ & _303_;
  assign _377_ = io_extendedMode & _321_;
  assign _379_ = _351_ & _378_;
  assign _380_ = _379_ & _357_;
  assign _382_ = _311_ & _381_;
  assign _383_ = io_extendedMode & _324_;
  assign _385_ = _351_ & _384_;
  assign _386_ = _385_ & _357_;
  assign read = io_cs & _310_;
  assign _388_ = _311_ & _387_;
  assign _390_ = _351_ & _389_;
  assign _391_ = _390_ & _357_;
  assign _393_ = _311_ & _392_;
  assign _394_ = io_extendedMode & _333_;
  assign _396_ = _351_ & _395_;
  assign _397_ = _396_ & _357_;
  assign _398_ = _311_ & _314_;
  assign _399_ = io_extendedMode & _336_;
  assign _401_ = _351_ & _400_;
  assign readIrqReg = read & _309_;
  assign _402_ = _401_ & _357_;
  assign _403_ = _311_ & _318_;
  assign _404_ = io_extendedMode & _339_;
  assign _406_ = _351_ & _405_;
  assign _407_ = _406_ & _357_;
  assign _408_ = _311_ & _321_;
  assign _410_ = io_extendedMode & _409_;
  assign _412_ = _351_ & _411_;
  assign _413_ = _412_ & _357_;
  assign _414_ = _311_ & _324_;
  assign _301_ = read & io_extendedMode;
  assign _416_ = io_extendedMode & _415_;
  assign _418_ = _351_ & _417_;
  assign _419_ = _418_ & _357_;
  assign _360_ = _351_ & _359_;
  assign _361_ = _360_ & io_extendedMode;
  assign _362_ = _361_ & _357_;
  assign _364_ = _351_ & _363_;
  assign _365_ = _364_ & io_extendedMode;
  assign _366_ = _365_ & _357_;
  assign _368_ = _351_ & _367_;
  assign _313_ = _311_ & _312_;
  assign _369_ = _368_ & io_extendedMode;
  assign _370_ = _369_ & _357_;
  assign _350_ = _351_ & _312_;
  assign _348_ = _351_ & _381_;
  assign _349_ = _348_ & io_extendedMode;
  assign _305_ = _351_ & _387_;
  assign _306_ = _305_ & io_extendedMode;
  assign _307_ = _351_ & _392_;
  assign _308_ = _307_ & io_extendedMode;
  assign _202_ = command_0 & io_samplePoint;
  assign _315_ = io_extendedMode & _314_;
  assign _204_ = io_abortTx & _203_;
  assign _206_ = io_samplePoint & _205_;
  assign _208_ = command_4 & io_samplePoint;
  assign _160_ = command_4 & _159_;
  assign _176_ = _170_ & io_txStateQ;
  assign _185_ = io_txRequest & command_1;
  assign _194_ = _185_ & io_samplePoint;
  assign _162_ = io_txSuccessful & _161_;
  assign _165_ = io_overrun & _164_;
  assign _171_ = _165_ & dataOverrunIrqEn;
  assign _317_ = _351_ & _316_;
  assign _174_ = transmitBufferStatus & _173_;
  assign _175_ = _174_ & transmitIrqEn;
  assign _178_ = _168_ & _177_;
  assign _179_ = _178_ & receiveIrqEn;
  assign _183_ = _182_ & errorWarningIrqEn;
  assign _184_ = io_setBusErrorIrq & busErrorIrqEn;
  assign _186_ = io_setArbitrationLostIrq & arbitrationLostIrqEn;
  assign _188_ = io_nodeErrorPassive & _187_;
  assign _190_ = _189_ & nodeErrorPassiveQ;
  assign _191_ = _190_ & io_nodeErrorActive;
  assign _352_ = ! io_addr;
  assign _347_ = io_addr == 8'h01;
  assign _342_ = io_addr == 8'h06;
  assign _329_ = io_addr == 8'h14;
  assign _318_ = io_addr == 8'h11;
  assign _333_ = io_addr == 8'h15;
  assign _321_ = io_addr == 8'h12;
  assign _336_ = io_addr == 8'h16;
  assign _324_ = io_addr == 8'h13;
  assign _339_ = io_addr == 8'h17;
  assign _353_ = io_addr == 8'h0a;
  assign _381_ = io_addr == 8'h0d;
  assign _387_ = io_addr == 8'h0e;
  assign _344_ = io_addr == 8'h07;
  assign _392_ = io_addr == 8'h0f;
  assign _409_ = io_addr == 8'h18;
  assign _415_ = io_addr == 8'h19;
  assign _359_ = io_addr == 8'h1a;
  assign _363_ = io_addr == 8'h1b;
  assign _367_ = io_addr == 8'h1c;
  assign _200_ = cd_m_io_dataOut == 3'h7;
  assign _169_ = clkoutCnt == clkoutDiv;
  assign _250_ = 5'h1f == _215_;
  assign _271_ = 5'h1d == _215_;
  assign _346_ = io_addr == 8'h1f;
  assign _284_ = 5'h17 == _215_;
  assign _217_ = 5'h16 == _215_;
  assign _220_ = 5'h15 == _215_;
  assign _222_ = 5'h14 == _215_;
  assign _224_ = 5'h13 == _215_;
  assign _226_ = 5'h12 == _215_;
  assign _229_ = 5'h11 == _215_;
  assign _231_ = 5'h10 == _215_;
  assign _233_ = 5'h0f == _215_;
  assign _235_ = 5'h0e == _215_;
  assign _309_ = io_addr == 8'h03;
  assign _237_ = 5'h0d == _215_;
  assign _240_ = 5'h0c == _215_;
  assign _242_ = 5'h0b == _215_;
  assign _244_ = 5'h07 == _215_;
  assign _246_ = 5'h06 == _215_;
  assign _248_ = 5'h04 == _215_;
  assign _251_ = 5'h03 == _215_;
  assign _253_ = 5'h02 == _215_;
  assign _255_ = ! _215_;
  assign _287_ = 5'h0a == _215_;
  assign _302_ = io_addr == 8'h0b;
  assign _292_ = 5'h05 == _215_;
  assign _297_ = 5'h01 == _215_;
  assign _303_ = io_addr == 8'h0c;
  assign _312_ = io_addr == 8'h04;
  assign _314_ = io_addr == 8'h10;
  assign _327_ = io_addr == 8'h05;
  assign _000_ = _176_ ? (* src = "CanRegisters.scala:182.43|CanRegisters.scala:183.19|CanRegisters.scala:102.36" *) 1'h0 : selfRxRequest;
  assign _011_ = _176_ ? (* src = "CanRegisters.scala:194.42|CanRegisters.scala:195.28|CanRegisters.scala:104.45" *) 1'h0 : singleShotTransmission;
  assign _025_ = io_txRequest ? (* src = "CanRegisters.scala:212.22|CanRegisters.scala:213.26" *) 1'h0 : _024_;
  assign _291_ = _284_ ? (* src = "Mux.scala:80.57" *) io_acceptanceMask_3 : _278_;
  assign _219_ = _217_ ? (* src = "Mux.scala:80.57" *) io_acceptanceMask_2 : _291_;
  assign _221_ = _220_ ? (* src = "Mux.scala:80.57" *) io_acceptanceMask_1 : _219_;
  assign _223_ = _222_ ? (* src = "Mux.scala:80.57" *) io_acceptanceMask_0 : _221_;
  assign _225_ = _224_ ? (* src = "Mux.scala:80.57" *) io_acceptanceCode_3 : _223_;
  assign _227_ = _226_ ? (* src = "Mux.scala:80.57" *) io_acceptanceCode_2 : _225_;
  assign _230_ = _229_ ? (* src = "Mux.scala:80.57" *) io_acceptanceCode_1 : _227_;
  assign _232_ = _231_ ? (* src = "Mux.scala:80.57" *) io_acceptanceCode_0 : _230_;
  assign _234_ = _233_ ? (* src = "Mux.scala:80.57" *) io_txErrorCount : _232_;
  assign _236_ = _235_ ? (* src = "Mux.scala:80.57" *) io_rxErrorCount : _234_;
  assign _026_ = io_txRequest ? (* src = "CanRegisters.scala:221.27|CanRegisters.scala:222.26|CanRegisters.scala:109.43" *) 1'h0 : transmissionComplete;
  assign _238_ = _237_ ? (* src = "Mux.scala:80.57" *) io_errorWarningLimit : _236_;
  assign _241_ = _240_ ? (* src = "Mux.scala:80.57" *) io_errorCaptureCode : _238_;
  assign _243_ = _242_ ? (* src = "Mux.scala:80.57" *) _228_ : _241_;
  assign _245_ = _244_ ? (* src = "Mux.scala:80.57" *) busTiming1_m_io_dataOut : _243_;
  assign _247_ = _246_ ? (* src = "Mux.scala:80.57" *) busTiming0_m_io_dataOut : _245_;
  assign _249_ = _248_ ? (* src = "Mux.scala:80.57" *) irqEnExt : _247_;
  assign _252_ = _251_ ? (* src = "Mux.scala:80.57" *) irqReg : _249_;
  assign _254_ = _253_ ? (* src = "Mux.scala:80.57" *) status : _252_;
  assign _256_ = _255_ ? (* src = "Mux.scala:80.57" *) _216_ : _254_;
  assign _261_ = io_resetMode ? (* src = "CanRegisters.scala:326.17" *) io_acceptanceCode_0 : 8'hff;
  assign _028_ = _166_ ? (* src = "CanRegisters.scala:228.49|CanRegisters.scala:229.19|CanRegisters.scala:108.36" *) 1'h0 : overrunStatus;
  assign _262_ = io_resetMode ? (* src = "CanRegisters.scala:327.17" *) io_acceptanceMask_0 : 8'hff;
  assign _263_ = io_resetMode ? (* src = "CanRegisters.scala:328.17" *) busTiming0_m_io_dataOut : 8'hff;
  assign _264_ = io_resetMode ? (* src = "CanRegisters.scala:329.17" *) busTiming1_m_io_dataOut : 8'hff;
  assign _265_ = io_resetMode ? (* src = "CanRegisters.scala:330.18" *) 8'hff : io_txData_0;
  assign _266_ = io_resetMode ? (* src = "CanRegisters.scala:331.18" *) 8'hff : io_txData_1;
  assign _267_ = io_resetMode ? (* src = "CanRegisters.scala:332.18" *) 8'hff : io_txData_2;
  assign _268_ = io_resetMode ? (* src = "CanRegisters.scala:333.18" *) 8'hff : io_txData_3;
  assign _269_ = io_resetMode ? (* src = "CanRegisters.scala:334.18" *) 8'hff : io_txData_4;
  assign _270_ = io_resetMode ? (* src = "CanRegisters.scala:335.18" *) 8'hff : io_txData_5;
  assign _272_ = io_resetMode ? (* src = "CanRegisters.scala:336.18" *) 8'hff : io_txData_6;
  assign _003_ = _167_ ? (* src = "CanRegisters.scala:232.41|CanRegisters.scala:233.25" *) 1'h0 : _002_;
  assign _273_ = io_resetMode ? (* src = "CanRegisters.scala:337.18" *) 8'hff : io_txData_7;
  assign _274_ = io_resetMode ? (* src = "CanRegisters.scala:338.18" *) 8'hff : io_txData_8;
  assign _275_ = io_resetMode ? (* src = "CanRegisters.scala:339.18" *) 8'hff : io_txData_9;
  assign _276_ = _224_ ? (* src = "Mux.scala:80.57" *) _275_ : _260_;
  assign _277_ = _226_ ? (* src = "Mux.scala:80.57" *) _274_ : _276_;
  assign _279_ = _229_ ? (* src = "Mux.scala:80.57" *) _273_ : _277_;
  assign _280_ = _231_ ? (* src = "Mux.scala:80.57" *) _272_ : _279_;
  assign _281_ = _233_ ? (* src = "Mux.scala:80.57" *) _270_ : _280_;
  assign _282_ = _235_ ? (* src = "Mux.scala:80.57" *) _269_ : _281_;
  assign _283_ = _237_ ? (* src = "Mux.scala:80.57" *) _268_ : _282_;
  assign clkoutDiv = _200_ ? (* src = "CanRegisters.scala:266.29" *) 3'h0 : cd_m_io_dataOut;
  assign _285_ = _240_ ? (* src = "Mux.scala:80.57" *) _267_ : _283_;
  assign _286_ = _242_ ? (* src = "Mux.scala:80.57" *) _266_ : _285_;
  assign _288_ = _287_ ? (* src = "Mux.scala:80.57" *) _265_ : _286_;
  assign _289_ = _244_ ? (* src = "Mux.scala:80.57" *) _264_ : _288_;
  assign _290_ = _246_ ? (* src = "Mux.scala:80.57" *) _263_ : _289_;
  assign _293_ = _292_ ? (* src = "Mux.scala:80.57" *) _262_ : _290_;
  assign _294_ = _248_ ? (* src = "Mux.scala:80.57" *) _261_ : _293_;
  assign _295_ = _251_ ? (* src = "Mux.scala:80.57" *) _259_ : _294_;
  assign _296_ = _253_ ? (* src = "Mux.scala:80.57" *) status : _295_;
  assign _298_ = _297_ ? (* src = "Mux.scala:80.57" *) 8'hff : _296_;
  assign _004_ = _169_ ? (* src = "CanRegisters.scala:271.33|CanRegisters.scala:272.15|CanRegisters.scala:276.15" *) 3'h0 : _199_;
  assign _218_ = _255_ ? (* src = "Mux.scala:80.57" *) _257_ : _298_;
  assign dataOverrunIrqEn = io_extendedMode ? (* src = "CanRegisters.scala:343.26" *) dataOverrunIrqEnExt : overrunIrqEnBasic;
  assign errorWarningIrqEn = io_extendedMode ? (* src = "CanRegisters.scala:344.27" *) errorWarningIrqEnExt : errorIrqEnBasic;
  assign transmitIrqEn = io_extendedMode ? (* src = "CanRegisters.scala:345.23" *) transmitIrqEnExt : transmitIrqEnBasic;
  assign receiveIrqEn = io_extendedMode ? (* src = "CanRegisters.scala:346.22" *) receiveIrqEnExt : receiveIrqEnBasic;
  assign _006_ = _172_ ? (* src = "CanRegisters.scala:358.41|CanRegisters.scala:359.20|CanRegisters.scala:348.38" *) 1'h0 : dataOverrunIrq;
  assign _009_ = _172_ ? (* src = "CanRegisters.scala:362.35|CanRegisters.scala:363.17" *) 1'h0 : _008_;
  assign _010_ = _167_ ? (* src = "CanRegisters.scala:370.48|CanRegisters.scala:371.16|CanRegisters.scala:350.34" *) 1'h0 : receiveIrq;
  assign _013_ = readIrqReg ? (* src = "CanRegisters.scala:376.26|CanRegisters.scala:377.14|CanRegisters.scala:351.32" *) 1'h0 : errorIrq;
  assign _015_ = _172_ ? (* src = "CanRegisters.scala:382.41|CanRegisters.scala:383.17|CanRegisters.scala:352.35" *) 1'h0 : busErrorIrq;
  assign _005_ = _169_ ? (* src = "CanRegisters.scala:271.33|CanRegisters.scala:273.15|CanRegisters.scala:269.33" *) _201_ : clkoutTmp;
  assign _017_ = _172_ ? (* src = "CanRegisters.scala:388.41|CanRegisters.scala:389.24|CanRegisters.scala:353.42" *) 1'h0 : arbitrationLostIrq;
  assign _019_ = _172_ ? (* src = "CanRegisters.scala:394.41|CanRegisters.scala:395.21|CanRegisters.scala:354.39" *) 1'h0 : errorPassiveIrq;
  assign _021_ = irq ? (* src = "CanRegisters.scala:403.19|CanRegisters.scala:404.10|CanRegisters.scala:100.27" *) 1'h0 : irqN;
  assign io_dataOut = io_extendedMode ? (* src = "CanRegisters.scala:297.20" *) _256_ : _218_;
  assign io_clkout = _211_ ? (* src = "CanRegisters.scala:281.31|CanRegisters.scala:282.16|CanRegisters.scala:285.15" *) _213_ : _214_;
  assign _260_ = _250_ ? (* src = "Mux.scala:80.57" *) clockDivider : 8'h00;
  assign _278_ = _271_ ? (* src = "Mux.scala:80.57" *) _239_ : _260_;
  assign _310_ = ~ io_writeEn;
  assign _311_ = ~ io_extendedMode;
  assign _357_ = ~ io_resetMode;
  assign _168_ = ~ io_infoEmpty;
  assign _201_ = ~ clkoutTmp;
  assign _173_ = ~ transmitBufferStatusQ;
  assign _177_ = ~ receiveIrq;
  assign _187_ = ~ nodeErrorPassiveQ;
  assign _189_ = ~ io_nodeErrorPassive;
  assign _203_ = ~ io_transmitting;
  assign _159_ = ~ command_0;
  assign _170_ = ~ io_txState;
  assign _209_ = ~ io_txRequest;
  assign _300_ = ~ overloadFrameQ;
  assign _196_ = ~ io_needToTx;
  assign _161_ = ~ txSuccessfulQ;
  assign _164_ = ~ overrunQ;
  assign _030_ = reset | _023_;
  assign _031_ = reset | _027_;
  assign _032_ = reset | _025_;
  assign _400_ = _398_ | _399_;
  assign _405_ = _403_ | _404_;
  assign _411_ = _408_ | _410_;
  assign _417_ = _414_ | _416_;
  assign _205_ = io_txRequest | _204_;
  assign _207_ = command_3 | command_2;
  assign _001_ = _160_ | _000_;
  assign _022_ = _194_ | _011_;
  assign _197_ = io_resetMode | _196_;
  assign _024_ = _197_ | transmitBufferStatus;
  assign _316_ = _313_ | _315_;
  assign _163_ = _162_ | io_abortTx;
  assign _027_ = _163_ | _026_;
  assign _166_ = io_resetMode | io_clearDataOverrun;
  assign _029_ = _165_ | _028_;
  assign _167_ = io_resetMode | io_releaseBuffer;
  assign _002_ = _168_ | receiveBufferStatus;
  assign _213_ = clockOff | _212_;
  assign _214_ = clockOff | clkoutTmp;
  assign _172_ = io_resetMode | readIrqReg;
  assign _007_ = _171_ | _006_;
  assign _331_ = _328_ | _330_;
  assign _008_ = _175_ | transmitIrq;
  assign _012_ = _179_ | _010_;
  assign _182_ = _180_ | _181_;
  assign _014_ = _183_ | _013_;
  assign _016_ = _184_ | _015_;
  assign _018_ = _186_ | _017_;
  assign _192_ = _188_ | _191_;
  assign _020_ = _193_ | _019_;
  assign _195_ = readIrqReg | io_releaseBuffer;
  assign _023_ = _195_ | _021_;
  assign _355_ = _354_ | _315_;
  assign io_txRequest = command_0 | command_4;
  assign _136_ = _202_ | io_resetMode;
  assign _140_ = _206_ | io_resetMode;
  assign _143_ = _207_ | io_resetMode;
  assign _146_ = _207_ | io_resetMode;
  assign _150_ = _208_ | io_resetMode;
  assign _373_ = _371_ | _372_;
  assign _378_ = _376_ | _377_;
  assign _384_ = _382_ | _383_;
  assign _389_ = _388_ | _330_;
  assign _395_ = _393_ | _394_;
  always @(posedge clock)
    receiveIrq <= _420_;
  always @(posedge clock)
    transmitIrq <= _422_;
  always @(posedge clock)
    errorIrq <= _424_;
  always @(posedge clock)
    dataOverrunIrq <= _426_;
  always @(posedge clock)
    errorPassiveIrq <= _428_;
  always @(posedge clock)
    arbitrationLostIrq <= _430_;
  always @(posedge clock)
    busErrorIrq <= _432_;
  always @(posedge clock)
    clkoutTmp <= _434_;
  always @(posedge clock)
    clkoutCnt <= _436_;
  always @(posedge clock)
    overloadFrameQ <= _438_;
  always @(posedge clock)
    nodeErrorPassiveQ <= io_nodeErrorPassive;
  always @(posedge clock)
    nodeBusOffQ <= io_nodeBusOff;
  always @(posedge clock)
    errorStatusQ <= io_errorStatus;
  always @(posedge clock)
    receiveBufferStatus <= _440_;
  always @(posedge clock)
    transmitBufferStatusQ <= transmitBufferStatus;
  always @(posedge clock)
    transmitBufferStatus <= _032_;
  always @(posedge clock)
    transmissionComplete <= _031_;
  always @(posedge clock)
    overrunStatus <= _442_;
  always @(posedge clock)
    overrunQ <= io_overrun;
  always @(posedge clock)
    txSuccessfulQ <= io_txSuccessful;
  always @(posedge clock)
    singleShotTransmission <= _444_;
  always @(posedge clock)
    selfRxRequest <= _446_;
  always @(posedge clock)
    irqN <= _030_;
  assign _420_ = _421_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:350.34" *) 1'h0 : _012_;
  assign _422_ = _423_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:349.35" *) 1'h0 : _009_;
  assign _424_ = _425_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:351.32" *) 1'h0 : _014_;
  assign _426_ = _427_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:348.38" *) 1'h0 : _007_;
  assign _428_ = _429_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:354.39" *) 1'h0 : _020_;
  assign _430_ = _431_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:353.42" *) 1'h0 : _018_;
  assign _432_ = _433_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:352.35" *) 1'h0 : _016_;
  assign _434_ = _435_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:269.33" *) 1'h0 : _005_;
  assign _436_ = _437_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:268.33" *) 3'h0 : _004_;
  assign _438_ = _439_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:198.38" *) 1'h0 : io_overloadFrame;
  assign _440_ = _441_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:112.42" *) 1'h0 : _003_;
  assign _442_ = _443_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:108.36" *) 1'h0 : _029_;
  assign _444_ = _445_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:104.45" *) 1'h0 : _022_;
  assign _446_ = _447_ ? (* full_case = 32'd1 *) (* src = "CanRegisters.scala:102.36" *) 1'h0 : _001_;
  assign _211_ = & cd_m_io_dataOut;
  assign irq = | irqReg;
  assign _180_ = io_errorStatus ^ errorStatusQ;
  assign _181_ = io_nodeBusOff ^ nodeBusOffQ;
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 busTiming0_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(busTiming0_m_io_dataOut),
    .io_writeEn(_157_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 busTiming1_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(busTiming1_m_io_dataOut),
    .io_writeEn(_158_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:30.19" *)
  CanRegister_1 cd_m (
    .clock(clock),
    .io_dataIn(io_dataIn[2:0]),
    .io_dataOut(cd_m_io_dataOut),
    .io_writeEn(_040_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:30.19" *)
  CanRegister_6 clockOff_m (
    .clock(clock),
    .io_dataIn(io_dataIn[3]),
    .io_dataOut(clockOff_m_io_dataOut),
    .io_writeEn(_038_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegisterDoubleReset.scala:24.19" *)
  CanRegisterDoubleReset_1 command_0_m (
    .clock(clock),
    .io_dataIn(io_dataIn[0]),
    .io_dataOut(command_0_m_io_dataOut),
    .io_resetSync(_136_),
    .io_writeEn(_139_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegisterDoubleReset.scala:24.19" *)
  CanRegisterDoubleReset_1 command_1_m (
    .clock(clock),
    .io_dataIn(io_dataIn[1]),
    .io_dataOut(command_1_m_io_dataOut),
    .io_resetSync(_140_),
    .io_writeEn(_142_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegisterDoubleReset.scala:24.19" *)
  CanRegisterDoubleReset_1 command_2_m (
    .clock(clock),
    .io_dataIn(io_dataIn[2]),
    .io_dataOut(command_2_m_io_dataOut),
    .io_resetSync(_143_),
    .io_writeEn(_145_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegisterDoubleReset.scala:24.19" *)
  CanRegisterDoubleReset_1 command_3_m (
    .clock(clock),
    .io_dataIn(io_dataIn[3]),
    .io_dataOut(command_3_m_io_dataOut),
    .io_resetSync(_146_),
    .io_writeEn(_149_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegisterDoubleReset.scala:24.19" *)
  CanRegisterDoubleReset_1 command_4_m (
    .clock(clock),
    .io_dataIn(io_dataIn[4]),
    .io_dataOut(command_4_m_io_dataOut),
    .io_resetSync(_150_),
    .io_writeEn(_152_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceCode_0_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceCode_0_m_io_dataOut),
    .io_writeEn(_041_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceCode_1_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceCode_1_m_io_dataOut),
    .io_writeEn(_043_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceCode_2_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceCode_2_m_io_dataOut),
    .io_writeEn(_046_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceCode_3_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceCode_3_m_io_dataOut),
    .io_writeEn(_048_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceMask_0_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceMask_0_m_io_dataOut),
    .io_writeEn(_042_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceMask_1_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceMask_1_m_io_dataOut),
    .io_writeEn(_045_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceMask_2_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceMask_2_m_io_dataOut),
    .io_writeEn(_047_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_acceptanceMask_3_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_acceptanceMask_3_m_io_dataOut),
    .io_writeEn(_049_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:30.19" *)
  CanRegister_5 io_errorWarningLimit_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_errorWarningLimit_m_io_dataOut),
    .io_writeEn(_034_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:30.19" *)
  CanRegister_6 io_extendedMode_m (
    .clock(clock),
    .io_dataIn(io_dataIn[7]),
    .io_dataOut(io_extendedMode_m_io_dataOut),
    .io_writeEn(_036_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegisterDoubleReset.scala:24.19" *)
  CanRegisterDoubleReset_1 io_overloadRequest_m (
    .clock(clock),
    .io_dataIn(io_dataIn[5]),
    .io_resetSync(_153_),
    .io_writeEn(_155_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_0_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_0_m_io_dataOut),
    .io_writeEn(_050_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_10_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_10_m_io_dataOut),
    .io_writeEn(_061_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_11_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_11_m_io_dataOut),
    .io_writeEn(_062_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_12_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_12_m_io_dataOut),
    .io_writeEn(_063_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_1_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_1_m_io_dataOut),
    .io_writeEn(_051_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_2_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_2_m_io_dataOut),
    .io_writeEn(_052_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_3_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_3_m_io_dataOut),
    .io_writeEn(_053_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_4_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_4_m_io_dataOut),
    .io_writeEn(_054_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_5_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_5_m_io_dataOut),
    .io_writeEn(_056_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_6_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_6_m_io_dataOut),
    .io_writeEn(_057_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_7_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_7_m_io_dataOut),
    .io_writeEn(_058_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_8_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_8_m_io_dataOut),
    .io_writeEn(_059_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 io_txData_9_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(io_txData_9_m_io_dataOut),
    .io_writeEn(_060_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:24.19" *)
  CanRegister_2 irqEnExt_m (
    .clock(clock),
    .io_dataIn(io_dataIn),
    .io_dataOut(irqEnExt_m_io_dataOut),
    .io_writeEn(_156_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:30.19" *)
  CanRegister modeBasic_m (
    .clock(clock),
    .io_dataIn(io_dataIn[4:1]),
    .io_dataOut(modeBasic_m_io_dataOut),
    .io_writeEn(_133_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegister.scala:30.19" *)
  CanRegister_1 modeExt_m (
    .clock(clock),
    .io_dataIn(io_dataIn[3:1]),
    .io_dataOut(modeExt_m_io_dataOut),
    .io_writeEn(_135_),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanRegisterDoubleReset.scala:24.19" *)
  CanRegisterDoubleReset mode_m (
    .clock(clock),
    .io_dataIn(io_dataIn[0]),
    .io_dataOut(mode_m_io_dataOut),
    .io_resetSync(io_setResetMode),
    .io_writeEn(_131_),
    .reset(reset)
  );
  assign mode = mode_m_io_dataOut;
  assign receiveIrqEnBasic = modeBasic_m_io_dataOut[0];
  assign transmitIrqEnBasic = modeBasic_m_io_dataOut[1];
  assign errorIrqEnBasic = modeBasic_m_io_dataOut[2];
  assign overrunIrqEnBasic = modeBasic_m_io_dataOut[3];
  assign _299_ = modeExt_m_io_dataOut[0];
  assign _304_ = modeExt_m_io_dataOut[1];
  assign _210_ = modeExt_m_io_dataOut[2];
  assign command_0 = command_0_m_io_dataOut;
  assign command_3 = command_3_m_io_dataOut;
  assign command_2 = command_2_m_io_dataOut;
  assign command_4 = command_4_m_io_dataOut;
  assign command_1 = command_1_m_io_dataOut;
  assign status = { io_nodeBusOff, io_errorStatus, io_transmitStatus, io_receiveStatus, transmissionComplete, transmitBufferStatus, overrunStatus, receiveBufferStatus };
  assign irqEnExt = irqEnExt_m_io_dataOut;
  assign busErrorIrqEn = irqEnExt[7];
  assign arbitrationLostIrqEn = irqEnExt[6];
  assign errorPassiveIrqEn = irqEnExt[5];
  assign dataOverrunIrqEnExt = irqEnExt[3];
  assign errorWarningIrqEnExt = irqEnExt[2];
  assign transmitIrqEnExt = irqEnExt[1];
  assign receiveIrqEnExt = irqEnExt[0];
  assign clockOff = clockOff_m_io_dataOut;
  assign clockDivider = { io_extendedMode, 3'h0, clockOff, cd_m_io_dataOut };
  assign _199_ = _198_[2:0];
  assign _212_ = clock;
  assign _215_ = io_addr[4:0];
  assign _216_ = { 4'h0, modeExt_m_io_dataOut, mode };
  assign _228_ = { 3'h0, io_arbitrationLostCapture };
  assign _239_ = { 1'h0, io_rxMessageCounter };
  assign irqReg = { busErrorIrq, arbitrationLostIrq, errorPassiveIrq, 1'h0, dataOverrunIrq, errorIrq, transmitIrq, receiveIrq };
  assign _257_ = { 3'h1, modeBasic_m_io_dataOut, mode };
  assign _258_ = irqReg[3:0];
  assign _259_ = { 4'he, _258_ };
  assign io_irqN = irqN;
  assign io_resetMode = mode_m_io_dataOut;
  assign io_clearDataOverrun = command_3_m_io_dataOut;
  assign io_releaseBuffer = command_2_m_io_dataOut;
  assign io_selfRxRequest = selfRxRequest;
  assign io_singleShotTransmission = singleShotTransmission;
  assign io_baudRatePrescaler = busTiming0_m_io_dataOut[5:0];
  assign io_syncJumpWidth = busTiming0_m_io_dataOut[7:6];
  assign io_timeSegment1 = busTiming1_m_io_dataOut[3:0];
  assign io_timeSegment2 = busTiming1_m_io_dataOut[6:4];
  assign io_tripleSampling = busTiming1_m_io_dataOut[7];
  assign io_errorWarningLimit = io_errorWarningLimit_m_io_dataOut;
  assign io_extendedMode = io_extendedMode_m_io_dataOut;
  assign io_acceptanceCode_0 = io_acceptanceCode_0_m_io_dataOut;
  assign io_acceptanceCode_1 = io_acceptanceCode_1_m_io_dataOut;
  assign io_acceptanceCode_2 = io_acceptanceCode_2_m_io_dataOut;
  assign io_acceptanceCode_3 = io_acceptanceCode_3_m_io_dataOut;
  assign io_acceptanceMask_0 = io_acceptanceMask_0_m_io_dataOut;
  assign io_acceptanceMask_1 = io_acceptanceMask_1_m_io_dataOut;
  assign io_acceptanceMask_2 = io_acceptanceMask_2_m_io_dataOut;
  assign io_acceptanceMask_3 = io_acceptanceMask_3_m_io_dataOut;
  assign io_txData_0 = io_txData_0_m_io_dataOut;
  assign io_txData_1 = io_txData_1_m_io_dataOut;
  assign io_txData_2 = io_txData_2_m_io_dataOut;
  assign io_txData_3 = io_txData_3_m_io_dataOut;
  assign io_txData_4 = io_txData_4_m_io_dataOut;
  assign io_txData_5 = io_txData_5_m_io_dataOut;
  assign io_txData_6 = io_txData_6_m_io_dataOut;
  assign io_txData_7 = io_txData_7_m_io_dataOut;
  assign io_txData_8 = io_txData_8_m_io_dataOut;
  assign io_txData_9 = io_txData_9_m_io_dataOut;
  assign io_txData_10 = io_txData_10_m_io_dataOut;
  assign io_txData_11 = io_txData_11_m_io_dataOut;
  assign io_txData_12 = io_txData_12_m_io_dataOut;
  assign \nodeErrorPassiveQ$process$CanRegisters_11  = io_nodeErrorPassive;
  assign \nodeBusOffQ$process$CanRegisters_10  = io_nodeBusOff;
  assign \errorStatusQ$process$CanRegisters_9  = io_errorStatus;
  assign \transmitBufferStatusQ$process$CanRegisters_7  = transmitBufferStatus;
  assign \transmitBufferStatus$process$CanRegisters_6  = _032_;
  assign \transmissionComplete$process$CanRegisters_5  = _031_;
  assign \overrunQ$process$CanRegisters_3  = io_overrun;
  assign \txSuccessfulQ$process$CanRegisters_2  = io_txSuccessful;
  assign \irqN$process$CanRegisters  = _030_;
  assign _421_ = reset;
  assign \receiveIrq$process$CanRegisters_21  = _420_;
  assign _423_ = reset;
  assign \transmitIrq$process$CanRegisters_20  = _422_;
  assign _425_ = reset;
  assign \errorIrq$process$CanRegisters_19  = _424_;
  assign _427_ = reset;
  assign \dataOverrunIrq$process$CanRegisters_18  = _426_;
  assign _429_ = reset;
  assign \errorPassiveIrq$process$CanRegisters_17  = _428_;
  assign _431_ = reset;
  assign \arbitrationLostIrq$process$CanRegisters_16  = _430_;
  assign _433_ = reset;
  assign \busErrorIrq$process$CanRegisters_15  = _432_;
  assign _435_ = reset;
  assign \clkoutTmp$process$CanRegisters_14  = _434_;
  assign _437_ = reset;
  assign \clkoutCnt$process$CanRegisters_13  = _436_;
  assign _439_ = reset;
  assign \overloadFrameQ$process$CanRegisters_12  = _438_;
  assign _441_ = reset;
  assign \receiveBufferStatus$process$CanRegisters_8  = _440_;
  assign _443_ = reset;
  assign \overrunStatus$process$CanRegisters_4  = _442_;
  assign _445_ = reset;
  assign \singleShotTransmission$process$CanRegisters_1  = _444_;
  assign _447_ = reset;
  assign \selfRxRequest$process$CanRegisters_0  = _446_;
endmodule

(* cells_not_processed =  1  *)
module CanTop(clock, reset, io_wbClkI, io_wbDatI, io_wbDatO, io_wbCycI, io_wbStbI, io_wbWeI, io_wbAddrI, io_wbAckO, io_canRx, io_canTx, io_busOffOn, io_irqOn, io_clkout);
  (* src = "CanTop.scala:285.19|CanTop.scala:286.10|CanTop.scala:95.28" *)
  wire [7:0] _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire [7:0] _04_;
  wire [7:0] _05_;
  (* src = "CanTop.scala:262.13" *)
  wire _06_;
  (* src = "CanTop.scala:262.11" *)
  wire _07_;
  (* src = "CanTop.scala:277.21" *)
  wire _08_;
  (* src = "CanTop.scala:276.25" *)
  wire _09_;
  (* src = "CanTop.scala:276.39" *)
  wire _10_;
  (* src = "CanTop.scala:276.37" *)
  wire _11_;
  (* src = "CanTop.scala:260.52" *)
  wire _12_;
  (* src = "CanTop.scala:260.49" *)
  wire _13_;
  (* src = "CanTop.scala:260.119" *)
  wire _14_;
  (* src = "CanTop.scala:260.73" *)
  wire _15_;
  (* src = "CanTop.scala:260.91" *)
  wire _16_;
  (* src = "CanTop.scala:260.82" *)
  wire _17_;
  (* src = "CanTop.scala:260.64" *)
  wire _18_;
  (* src = "CanTop.scala:260.104" *)
  wire _19_;
  (* src = "CanTop.scala:260.128" *)
  wire _20_;
  (* src = "CanTop.scala:260.146" *)
  wire _21_;
  (* src = "CanTop.scala:260.137" *)
  wire _22_;
  (* src = "CanTop.scala:263.21" *)
  wire [7:0] _23_;
  (* src = "CanTop.scala:280.24" *)
  wire _24_;
  (* src = "CanTop.scala:280.21" *)
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire [7:0] _38_;
  wire _39_;
  wire _40_;
  wire [7:0] _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  (* src = "CanTop.scala:95.28" *)
  reg [7:0] addr;
  (* src = "CanTop.scala:95.28|CanTop.scala:95.28" *)
  wire [7:0] \addr$process$CanTop ;
  (* src = "CanTop.scala:84.43|CanTop.scala:240.26" *)
  wire [4:0] canBsp_io_arbitrationLostCapture;
  (* src = "CanTop.scala:246.15" *)
  wire canBsp_io_busOffOn;
  (* src = "CanTop.scala:21.32|CanTop.scala:197.15" *)
  wire [7:0] canBsp_io_dataOut;
  (* src = "CanTop.scala:41.37|CanTop.scala:215.20" *)
  wire [7:0] canBsp_io_errorCaptureCode;
  (* src = "CanTop.scala:73.31|CanTop.scala:229.15" *)
  wire canBsp_io_errorStatus;
  (* src = "CanTop.scala:91.33|CanTop.scala:248.16" *)
  wire canBsp_io_goErrorFrame;
  (* src = "CanTop.scala:90.36|CanTop.scala:247.19" *)
  wire canBsp_io_goOverloadFrame;
  (* src = "CanTop.scala:68.30|CanTop.scala:224.13" *)
  wire canBsp_io_goRxInter;
  (* src = "CanTop.scala:92.25|CanTop.scala:249.8" *)
  wire canBsp_io_goTx;
  (* src = "CanTop.scala:81.30|CanTop.scala:237.13" *)
  wire canBsp_io_infoEmpty;
  (* src = "CanTop.scala:79.29|CanTop.scala:235.12" *)
  wire canBsp_io_needToTx;
  (* src = "CanTop.scala:72.31|CanTop.scala:228.14" *)
  wire canBsp_io_nodeBusOff;
  (* src = "CanTop.scala:86.36|CanTop.scala:242.19" *)
  wire canBsp_io_nodeErrorActive;
  (* src = "CanTop.scala:85.37|CanTop.scala:241.20" *)
  wire canBsp_io_nodeErrorPassive;
  (* src = "CanTop.scala:36.34|CanTop.scala:210.17" *)
  wire canBsp_io_overloadFrame;
  (* src = "CanTop.scala:80.28|CanTop.scala:236.11" *)
  wire canBsp_io_overrun;
  (* src = "CanTop.scala:77.34|CanTop.scala:233.17" *)
  wire canBsp_io_receiveStatus;
  wire [8:0] canBsp_io_rxErrorCount;
  (* src = "CanTop.scala:65.27|CanTop.scala:222.10" *)
  wire canBsp_io_rxIdle;
  (* src = "CanTop.scala:69.28|CanTop.scala:226.11" *)
  wire canBsp_io_rxInter;
  (* src = "CanTop.scala:87.37|CanTop.scala:243.20" *)
  wire [6:0] canBsp_io_rxMessageCounter;
  (* src = "CanTop.scala:93.28|CanTop.scala:250.11" *)
  wire canBsp_io_sendAck;
  (* src = "CanTop.scala:83.42|CanTop.scala:239.25" *)
  wire canBsp_io_setArbitrationLostIrq;
  (* src = "CanTop.scala:82.35|CanTop.scala:238.18" *)
  wire canBsp_io_setBusErrorIrq;
  (* src = "CanTop.scala:71.33|CanTop.scala:227.16" *)
  wire canBsp_io_setResetMode;
  (* src = "CanTop.scala:76.35|CanTop.scala:232.18" *)
  wire canBsp_io_transmitStatus;
  (* src = "CanTop.scala:67.32|CanTop.scala:251.15" *)
  wire canBsp_io_transmitter;
  (* src = "CanTop.scala:66.33|CanTop.scala:252.16" *)
  wire canBsp_io_transmitting;
  (* src = "CanTop.scala:244.12" *)
  wire canBsp_io_tx;
  wire [8:0] canBsp_io_txErrorCount;
  (* src = "CanTop.scala:88.27|CanTop.scala:245.10" *)
  wire canBsp_io_txNext;
  (* src = "CanTop.scala:34.28|CanTop.scala:207.11" *)
  wire canBsp_io_txState;
  (* src = "CanTop.scala:35.29|CanTop.scala:208.12" *)
  wire canBsp_io_txStateQ;
  (* src = "CanTop.scala:78.33|CanTop.scala:253.16" *)
  wire canBsp_io_txSuccessful;
  (* src = "CanTop.scala:194.22" *)
  wire canBtl_io_hardSync;
  (* src = "CanTop.scala:59.32|CanTop.scala:171.15" *)
  wire canBtl_io_samplePoint;
  (* src = "CanTop.scala:191.24" *)
  wire canBtl_io_sampledBit;
  (* src = "CanTop.scala:192.25" *)
  wire canBtl_io_sampledBitQ;
  (* src = "CanTop.scala:193.21" *)
  wire canBtl_io_txPoint;
  (* src = "CanTop.scala:203.21" *)
  wire canRegisters_io_abortTx;
  (* src = "CanTop.scala:255.28" *)
  wire [7:0] canRegisters_io_acceptanceCode_0;
  (* src = "CanTop.scala:255.28" *)
  wire [7:0] canRegisters_io_acceptanceCode_1;
  (* src = "CanTop.scala:255.28" *)
  wire [7:0] canRegisters_io_acceptanceCode_2;
  (* src = "CanTop.scala:255.28" *)
  wire [7:0] canRegisters_io_acceptanceCode_3;
  (* src = "CanTop.scala:26.41|CanTop.scala:129.24" *)
  wire canRegisters_io_acceptanceFilterMode;
  (* src = "CanTop.scala:256.28" *)
  wire [7:0] canRegisters_io_acceptanceMask_0;
  (* src = "CanTop.scala:256.28" *)
  wire [7:0] canRegisters_io_acceptanceMask_1;
  (* src = "CanTop.scala:256.28" *)
  wire [7:0] canRegisters_io_acceptanceMask_2;
  (* src = "CanTop.scala:256.28" *)
  wire [7:0] canRegisters_io_acceptanceMask_3;
  (* src = "CanTop.scala:43.38|CanTop.scala:146.21" *)
  wire [5:0] canRegisters_io_baudRatePrescaler;
  (* src = "CanTop.scala:158.13" *)
  wire canRegisters_io_clkout;
  (* src = "CanTop.scala:22.32|CanTop.scala:106.15" *)
  wire [7:0] canRegisters_io_dataOut;
  (* src = "CanTop.scala:49.38|CanTop.scala:153.21" *)
  wire [7:0] canRegisters_io_errorWarningLimit;
  (* src = "CanTop.scala:55.33|CanTop.scala:157.16" *)
  wire canRegisters_io_extendedMode;
  (* src = "CanTop.scala:107.12" *)
  wire canRegisters_io_irqN;
  (* src = "CanTop.scala:25.35|CanTop.scala:128.18" *)
  wire canRegisters_io_listenOnlyMode;
  (* src = "CanTop.scala:212.43" *)
  wire canRegisters_io_readArbitrationLostCaptureReg;
  (* src = "CanTop.scala:214.37" *)
  wire canRegisters_io_readErrorCodeCaptureReg;
  (* src = "CanTop.scala:202.27" *)
  wire canRegisters_io_releaseBuffer;
  (* src = "CanTop.scala:24.30|CanTop.scala:127.13" *)
  wire canRegisters_io_resetMode;
  (* src = "CanTop.scala:205.27" *)
  wire canRegisters_io_selfRxRequest;
  (* src = "CanTop.scala:27.33|CanTop.scala:130.16" *)
  wire canRegisters_io_selfTestMode;
  (* src = "CanTop.scala:206.36" *)
  wire canRegisters_io_singleShotTransmission;
  (* src = "CanTop.scala:44.34|CanTop.scala:147.17" *)
  wire [1:0] canRegisters_io_syncJumpWidth;
  (* src = "CanTop.scala:45.33|CanTop.scala:149.16" *)
  wire [3:0] canRegisters_io_timeSegment1;
  (* src = "CanTop.scala:46.33|CanTop.scala:150.16" *)
  wire [2:0] canRegisters_io_timeSegment2;
  (* src = "CanTop.scala:47.35|CanTop.scala:151.18" *)
  wire canRegisters_io_tripleSampling;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_0;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_1;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_10;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_11;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_12;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_2;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_3;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_4;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_5;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_6;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_7;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_8;
  (* src = "CanTop.scala:258.20" *)
  wire [7:0] canRegisters_io_txData_9;
  (* src = "CanTop.scala:204.23" *)
  wire canRegisters_io_txRequest;
  (* src = "CanTop.scala:218.40" *)
  wire canRegisters_io_writeEnReceiveErrorCounter;
  (* src = "CanTop.scala:219.41" *)
  wire canRegisters_io_writeEnTransmitErrorCounter;
  input clock;
  (* src = "CanTop.scala:277.18" *)
  wire cs;
  (* src = "CanTop.scala:270.53" *)
  reg cs_ack1;
  (* src = "CanTop.scala:270.53|CanTop.scala:270.53|CanTop.scala:270.53" *)
  wire \cs_ack1$process$CanTop_6 ;
  (* src = "CanTop.scala:271.53" *)
  reg cs_ack2;
  (* src = "CanTop.scala:271.53|CanTop.scala:271.53|CanTop.scala:271.53" *)
  wire \cs_ack2$process$CanTop_7 ;
  (* src = "CanTop.scala:272.53" *)
  reg cs_ack3;
  (* src = "CanTop.scala:272.53|CanTop.scala:272.53|CanTop.scala:272.53" *)
  wire \cs_ack3$process$CanTop_8 ;
  (* src = "CanTop.scala:266.31" *)
  reg cs_sync1;
  (* src = "CanTop.scala:266.31|CanTop.scala:266.31|CanTop.scala:276.12" *)
  wire \cs_sync1$process$CanTop_5 ;
  (* src = "CanTop.scala:267.31" *)
  reg cs_sync2;
  (* src = "CanTop.scala:267.31|CanTop.scala:267.31|CanTop.scala:267.31" *)
  wire \cs_sync2$process$CanTop_3 ;
  (* src = "CanTop.scala:268.31" *)
  reg cs_sync3;
  (* src = "CanTop.scala:268.31|CanTop.scala:268.31|CanTop.scala:268.31" *)
  wire \cs_sync3$process$CanTop_4 ;
  (* src = "CanTop.scala:274.35" *)
  reg cs_sync_rst1;
  (* src = "CanTop.scala:274.35|CanTop.scala:274.35|CanTop.scala:274.35" *)
  wire \cs_sync_rst1$process$CanTop_9 ;
  (* src = "CanTop.scala:275.35" *)
  reg cs_sync_rst2;
  (* src = "CanTop.scala:275.35|CanTop.scala:275.35|CanTop.scala:275.35" *)
  wire \cs_sync_rst2$process$CanTop_10 ;
  (* src = "CanTop.scala:97.27" *)
  reg [7:0] dataOut;
  (* src = "CanTop.scala:262.23|CanTop.scala:263.15|CanTop.scala:97.27" *)
  wire [7:0] \dataOut$process$CanTop_0 ;
  (* src = "CanTop.scala:21.32|CanTop.scala:197.15" *)
  wire [7:0] dataOutFifo;
  (* src = "CanTop.scala:260.101" *)
  wire dataOutFifoSelected;
  (* src = "CanTop.scala:22.32|CanTop.scala:106.15" *)
  wire [7:0] dataOutRegs;
  (* src = "CanTop.scala:55.33|CanTop.scala:157.16" *)
  wire extendedMode;
  output io_busOffOn;
  input io_canRx;
  output io_canTx;
  output io_clkout;
  output io_irqOn;
  output io_wbAckO;
  input [7:0] io_wbAddrI;
  input io_wbClkI;
  input io_wbCycI;
  input [7:0] io_wbDatI;
  output [7:0] io_wbDatO;
  input io_wbStbI;
  input io_wbWeI;
  input reset;
  (* src = "CanTop.scala:24.30|CanTop.scala:127.13" *)
  wire resetMode;
  (* src = "CanTop.scala:99.30" *)
  reg rxSync;
  (* src = "CanTop.scala:99.30|CanTop.scala:99.30|CanTop.scala:99.30" *)
  wire \rxSync$process$CanTop_2 ;
  (* src = "CanTop.scala:98.33" *)
  reg rxSyncTmp;
  (* src = "CanTop.scala:98.33|CanTop.scala:98.33|CanTop.scala:98.33" *)
  wire \rxSyncTmp$process$CanTop_1 ;
  (* src = "CanTop.scala:280.12" *)
  reg wbAckO;
  (* src = "CanTop.scala:280.12|CanTop.scala:280.12|CanTop.scala:280.12" *)
  wire \wbAckO$process$CanTop_11 ;
  assign _13_ = extendedMode & _12_;
  assign _17_ = _15_ & _16_;
  assign _18_ = _13_ & _17_;
  assign _22_ = _20_ & _21_;
  assign _14_ = _19_ & _22_;
  assign cs = cs_sync2 & _08_;
  assign _07_ = cs & _06_;
  assign _09_ = io_wbCycI & io_wbStbI;
  assign _11_ = _09_ & _10_;
  assign _25_ = cs_ack2 & _24_;
  assign _03_ = cs_sync2 & _08_;
  assign _15_ = addr >= 8'h10;
  assign _20_ = addr >= 8'h14;
  assign _16_ = addr <= 8'h1c;
  assign _21_ = addr <= 8'h1d;
  assign _23_ = dataOutFifoSelected ? (* src = "CanTop.scala:263.21" *) dataOutFifo : dataOutRegs;
  assign _00_ = io_wbStbI ? (* src = "CanTop.scala:285.19|CanTop.scala:286.10|CanTop.scala:95.28" *) io_wbAddrI : addr;
  assign _12_ = ~ resetMode;
  assign _19_ = ~ extendedMode;
  assign _06_ = ~ io_wbWeI;
  assign _08_ = ~ cs_sync3;
  assign _10_ = ~ cs_sync_rst2;
  assign _24_ = ~ cs_ack3;
  assign _01_ = reset | io_canRx;
  assign _02_ = reset | rxSyncTmp;
  assign dataOutFifoSelected = _18_ | _14_;
  always @(posedge io_wbClkI)
    wbAckO <= _40_;
  always @(posedge clock)
    cs_sync_rst2 <= _44_;
  always @(posedge clock)
    cs_sync_rst1 <= _46_;
  always @(posedge io_wbClkI)
    cs_ack3 <= _26_;
  always @(posedge io_wbClkI)
    cs_ack2 <= _28_;
  always @(posedge io_wbClkI)
    cs_ack1 <= _30_;
  always @(posedge clock)
    cs_sync1 <= _32_;
  always @(posedge clock)
    cs_sync3 <= _34_;
  always @(posedge clock)
    cs_sync2 <= _36_;
  always @(posedge clock)
    rxSync <= _02_;
  always @(posedge clock)
    rxSyncTmp <= _01_;
  always @(posedge clock)
    dataOut <= _38_;
  always @(posedge clock)
    addr <= _41_;
  assign _26_ = _27_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:272.53" *) 1'h0 : cs_ack2;
  assign _28_ = _29_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:271.53" *) 1'h0 : cs_ack1;
  assign _30_ = _31_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:270.53" *) 1'h0 : cs_sync3;
  assign _40_ = _43_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:280.12" *) 1'h0 : _25_;
  assign _32_ = _33_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:266.31" *) 1'h0 : _11_;
  assign _34_ = _35_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:268.31" *) 1'h0 : cs_sync2;
  assign _36_ = _37_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:267.31" *) 1'h0 : cs_sync1;
  assign _38_ = _39_ ? (* src = "CanTop.scala:263.15|CanTop.scala:262.23" *) _23_ : dataOut;
  assign _41_ = _42_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:95.28" *) 8'h00 : _00_;
  assign _44_ = _45_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:275.35" *) 1'h0 : cs_sync_rst1;
  assign _46_ = _47_ ? (* full_case = 32'd1 *) (* src = "CanTop.scala:274.35" *) 1'h0 : cs_ack3;
  (* module_not_derived = 32'd1 *)
  (* src = "CanTop.scala:189.31" *)
  CanBsp canBsp (
    .clock(clock),
    .io_abortTx(canRegisters_io_abortTx),
    .io_acceptanceCode_0(canRegisters_io_acceptanceCode_0),
    .io_acceptanceCode_1(canRegisters_io_acceptanceCode_1),
    .io_acceptanceCode_2(canRegisters_io_acceptanceCode_2),
    .io_acceptanceCode_3(canRegisters_io_acceptanceCode_3),
    .io_acceptanceFilterMode(canRegisters_io_acceptanceFilterMode),
    .io_acceptanceMask_0(canRegisters_io_acceptanceMask_0),
    .io_acceptanceMask_1(canRegisters_io_acceptanceMask_1),
    .io_acceptanceMask_2(canRegisters_io_acceptanceMask_2),
    .io_acceptanceMask_3(canRegisters_io_acceptanceMask_3),
    .io_addr(addr),
    .io_arbitrationLostCapture(canBsp_io_arbitrationLostCapture),
    .io_busOffOn(canBsp_io_busOffOn),
    .io_dataIn(io_wbDatI),
    .io_dataOut(canBsp_io_dataOut),
    .io_errorCaptureCode(canBsp_io_errorCaptureCode),
    .io_errorStatus(canBsp_io_errorStatus),
    .io_errorWarningLimit(canRegisters_io_errorWarningLimit),
    .io_extendedMode(canRegisters_io_extendedMode),
    .io_goErrorFrame(canBsp_io_goErrorFrame),
    .io_goOverloadFrame(canBsp_io_goOverloadFrame),
    .io_goRxInter(canBsp_io_goRxInter),
    .io_goTx(canBsp_io_goTx),
    .io_hardSync(canBtl_io_hardSync),
    .io_infoEmpty(canBsp_io_infoEmpty),
    .io_listenOnlyMode(canRegisters_io_listenOnlyMode),
    .io_needToTx(canBsp_io_needToTx),
    .io_nodeBusOff(canBsp_io_nodeBusOff),
    .io_nodeErrorActive(canBsp_io_nodeErrorActive),
    .io_nodeErrorPassive(canBsp_io_nodeErrorPassive),
    .io_overloadFrame(canBsp_io_overloadFrame),
    .io_overrun(canBsp_io_overrun),
    .io_readArbitrationLostCaptureReg(canRegisters_io_readArbitrationLostCaptureReg),
    .io_readErrorCodeCaptureReg(canRegisters_io_readErrorCodeCaptureReg),
    .io_receiveStatus(canBsp_io_receiveStatus),
    .io_releaseBuffer(canRegisters_io_releaseBuffer),
    .io_resetMode(canRegisters_io_resetMode),
    .io_rxErrorCount(canBsp_io_rxErrorCount),
    .io_rxIdle(canBsp_io_rxIdle),
    .io_rxInter(canBsp_io_rxInter),
    .io_rxMessageCounter(canBsp_io_rxMessageCounter),
    .io_samplePoint(canBtl_io_samplePoint),
    .io_sampledBit(canBtl_io_sampledBit),
    .io_sampledBitQ(canBtl_io_sampledBitQ),
    .io_selfRxRequest(canRegisters_io_selfRxRequest),
    .io_selfTestMode(canRegisters_io_selfTestMode),
    .io_sendAck(canBsp_io_sendAck),
    .io_setArbitrationLostIrq(canBsp_io_setArbitrationLostIrq),
    .io_setBusErrorIrq(canBsp_io_setBusErrorIrq),
    .io_setResetMode(canBsp_io_setResetMode),
    .io_singleShotTransmission(canRegisters_io_singleShotTransmission),
    .io_transmitStatus(canBsp_io_transmitStatus),
    .io_transmitter(canBsp_io_transmitter),
    .io_transmitting(canBsp_io_transmitting),
    .io_tx(canBsp_io_tx),
    .io_txData_0(canRegisters_io_txData_0),
    .io_txData_1(canRegisters_io_txData_1),
    .io_txData_10(canRegisters_io_txData_10),
    .io_txData_11(canRegisters_io_txData_11),
    .io_txData_12(canRegisters_io_txData_12),
    .io_txData_2(canRegisters_io_txData_2),
    .io_txData_3(canRegisters_io_txData_3),
    .io_txData_4(canRegisters_io_txData_4),
    .io_txData_5(canRegisters_io_txData_5),
    .io_txData_6(canRegisters_io_txData_6),
    .io_txData_7(canRegisters_io_txData_7),
    .io_txData_8(canRegisters_io_txData_8),
    .io_txData_9(canRegisters_io_txData_9),
    .io_txErrorCount(canBsp_io_txErrorCount),
    .io_txNext(canBsp_io_txNext),
    .io_txPoint(canBtl_io_txPoint),
    .io_txRequest(canRegisters_io_txRequest),
    .io_txState(canBsp_io_txState),
    .io_txStateQ(canBsp_io_txStateQ),
    .io_txSuccessful(canBsp_io_txSuccessful),
    .io_writeEnReceiveErrorCounter(canRegisters_io_writeEnReceiveErrorCounter),
    .io_writeEnTransmitErrorCounter(canRegisters_io_writeEnTransmitErrorCounter),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanTop.scala:160.31" *)
  CanBtl canBtl (
    .clock(clock),
    .io_baudRatePrescaler(canRegisters_io_baudRatePrescaler),
    .io_goErrorFrame(canBsp_io_goErrorFrame),
    .io_goOverloadFrame(canBsp_io_goOverloadFrame),
    .io_goRxInter(canBsp_io_goRxInter),
    .io_goTx(canBsp_io_goTx),
    .io_hardSync(canBtl_io_hardSync),
    .io_nodeErrorPassive(canBsp_io_nodeErrorPassive),
    .io_rx(rxSync),
    .io_rxIdle(canBsp_io_rxIdle),
    .io_rxInter(canBsp_io_rxInter),
    .io_samplePoint(canBtl_io_samplePoint),
    .io_sampledBit(canBtl_io_sampledBit),
    .io_sampledBitQ(canBtl_io_sampledBitQ),
    .io_sendAck(canBsp_io_sendAck),
    .io_syncJumpWidth(canRegisters_io_syncJumpWidth),
    .io_timeSegment1(canRegisters_io_timeSegment1),
    .io_timeSegment2(canRegisters_io_timeSegment2),
    .io_transmitter(canBsp_io_transmitter),
    .io_transmitting(canBsp_io_transmitting),
    .io_tripleSampling(canRegisters_io_tripleSampling),
    .io_tx(io_canTx),
    .io_txNext(canBsp_io_txNext),
    .io_txPoint(canBtl_io_txPoint),
    .reset(reset)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "CanTop.scala:101.43" *)
  CanRegisters canRegisters (
    .clock(clock),
    .io_abortTx(canRegisters_io_abortTx),
    .io_acceptanceCode_0(canRegisters_io_acceptanceCode_0),
    .io_acceptanceCode_1(canRegisters_io_acceptanceCode_1),
    .io_acceptanceCode_2(canRegisters_io_acceptanceCode_2),
    .io_acceptanceCode_3(canRegisters_io_acceptanceCode_3),
    .io_acceptanceFilterMode(canRegisters_io_acceptanceFilterMode),
    .io_acceptanceMask_0(canRegisters_io_acceptanceMask_0),
    .io_acceptanceMask_1(canRegisters_io_acceptanceMask_1),
    .io_acceptanceMask_2(canRegisters_io_acceptanceMask_2),
    .io_acceptanceMask_3(canRegisters_io_acceptanceMask_3),
    .io_addr(addr),
    .io_arbitrationLostCapture(canBsp_io_arbitrationLostCapture),
    .io_baudRatePrescaler(canRegisters_io_baudRatePrescaler),
    .io_clkout(canRegisters_io_clkout),
    .io_cs(_03_),
    .io_dataIn(io_wbDatI),
    .io_dataOut(canRegisters_io_dataOut),
    .io_errorCaptureCode(canBsp_io_errorCaptureCode),
    .io_errorStatus(canBsp_io_errorStatus),
    .io_errorWarningLimit(canRegisters_io_errorWarningLimit),
    .io_extendedMode(canRegisters_io_extendedMode),
    .io_infoEmpty(canBsp_io_infoEmpty),
    .io_irqN(canRegisters_io_irqN),
    .io_listenOnlyMode(canRegisters_io_listenOnlyMode),
    .io_needToTx(canBsp_io_needToTx),
    .io_nodeBusOff(canBsp_io_nodeBusOff),
    .io_nodeErrorActive(canBsp_io_nodeErrorActive),
    .io_nodeErrorPassive(canBsp_io_nodeErrorPassive),
    .io_overloadFrame(canBsp_io_overloadFrame),
    .io_overrun(canBsp_io_overrun),
    .io_readArbitrationLostCaptureReg(canRegisters_io_readArbitrationLostCaptureReg),
    .io_readErrorCodeCaptureReg(canRegisters_io_readErrorCodeCaptureReg),
    .io_receiveStatus(canBsp_io_receiveStatus),
    .io_releaseBuffer(canRegisters_io_releaseBuffer),
    .io_resetMode(canRegisters_io_resetMode),
    .io_rxErrorCount(canBsp_io_rxErrorCount[7:0]),
    .io_rxMessageCounter(canBsp_io_rxMessageCounter),
    .io_samplePoint(canBtl_io_samplePoint),
    .io_selfRxRequest(canRegisters_io_selfRxRequest),
    .io_selfTestMode(canRegisters_io_selfTestMode),
    .io_setArbitrationLostIrq(canBsp_io_setArbitrationLostIrq),
    .io_setBusErrorIrq(canBsp_io_setBusErrorIrq),
    .io_setResetMode(canBsp_io_setResetMode),
    .io_singleShotTransmission(canRegisters_io_singleShotTransmission),
    .io_syncJumpWidth(canRegisters_io_syncJumpWidth),
    .io_timeSegment1(canRegisters_io_timeSegment1),
    .io_timeSegment2(canRegisters_io_timeSegment2),
    .io_transmitStatus(canBsp_io_transmitStatus),
    .io_transmitting(canBsp_io_transmitting),
    .io_tripleSampling(canRegisters_io_tripleSampling),
    .io_txData_0(canRegisters_io_txData_0),
    .io_txData_1(canRegisters_io_txData_1),
    .io_txData_10(canRegisters_io_txData_10),
    .io_txData_11(canRegisters_io_txData_11),
    .io_txData_12(canRegisters_io_txData_12),
    .io_txData_2(canRegisters_io_txData_2),
    .io_txData_3(canRegisters_io_txData_3),
    .io_txData_4(canRegisters_io_txData_4),
    .io_txData_5(canRegisters_io_txData_5),
    .io_txData_6(canRegisters_io_txData_6),
    .io_txData_7(canRegisters_io_txData_7),
    .io_txData_8(canRegisters_io_txData_8),
    .io_txData_9(canRegisters_io_txData_9),
    .io_txErrorCount(canBsp_io_txErrorCount[7:0]),
    .io_txRequest(canRegisters_io_txRequest),
    .io_txState(canBsp_io_txState),
    .io_txStateQ(canBsp_io_txStateQ),
    .io_txSuccessful(canBsp_io_txSuccessful),
    .io_writeEn(io_wbWeI),
    .io_writeEnReceiveErrorCounter(canRegisters_io_writeEnReceiveErrorCounter),
    .io_writeEnTransmitErrorCounter(canRegisters_io_writeEnTransmitErrorCounter),
    .reset(reset)
  );
  assign resetMode = canRegisters_io_resetMode;
  assign extendedMode = canRegisters_io_extendedMode;
  assign dataOutFifo = canBsp_io_dataOut;
  assign dataOutRegs = canRegisters_io_dataOut;
  assign io_wbDatO = dataOut;
  assign io_wbAckO = wbAckO;
  assign io_canTx = canBsp_io_tx;
  assign io_busOffOn = canBsp_io_busOffOn;
  assign io_irqOn = canRegisters_io_irqN;
  assign io_clkout = canRegisters_io_clkout;
  assign \rxSync$process$CanTop_2  = _02_;
  assign \rxSyncTmp$process$CanTop_1  = _01_;
  assign _43_ = reset;
  assign \wbAckO$process$CanTop_11  = _40_;
  assign _45_ = reset;
  assign \cs_sync_rst2$process$CanTop_10  = _44_;
  assign _47_ = reset;
  assign \cs_sync_rst1$process$CanTop_9  = _46_;
  assign _27_ = reset;
  assign \cs_ack3$process$CanTop_8  = _26_;
  assign _29_ = reset;
  assign \cs_ack2$process$CanTop_7  = _28_;
  assign _31_ = reset;
  assign \cs_ack1$process$CanTop_6  = _30_;
  assign _33_ = reset;
  assign \cs_sync1$process$CanTop_5  = _32_;
  assign _35_ = reset;
  assign \cs_sync3$process$CanTop_4  = _34_;
  assign _37_ = reset;
  assign \cs_sync2$process$CanTop_3  = _36_;
  assign _39_ = _07_;
  assign \dataOut$process$CanTop_0  = _38_;
  assign _42_ = reset;
  assign \addr$process$CanTop  = _41_;
endmodule
`default_nettype none
